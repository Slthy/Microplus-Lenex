<?xml version="1.0" encoding="utf-8" standalone="no"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="Swiss Timing Swimming Data Handling" version="60.0.0.0">
    <CONTACT name="Swiss Timing Ltd." zip="CH-2606" city="Corgemont" email="info@swisstiming.com" internet="http://www.swisstiming.com" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET name="16th FINA World Swimming Championships (25m)" city="Melbourne" nation="AUS" course="SCM" timing="AUTOMATIC">
      <POOL lanemin="0" lanemax="10" />
      <POINTTABLE name="FINA Point Scoring" version="2004" />
      <SESSIONS>
        <SESSION number="1" date="2022-12-13" daytime="11:05">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="1" number="1" preveventid="-1" gender="F" round="PRE" daytime="11:05">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="11:06" heatid="10001" number="1" />
                <HEAT daytime="11:12" heatid="20001" number="2" />
                <HEAT daytime="11:18" heatid="30001" number="3" />
                <HEAT daytime="11:24" heatid="40001" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2" number="2" preveventid="-1" gender="F" round="PRE" daytime="11:28">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="11:41" heatid="10002" number="1" />
                <HEAT daytime="11:44" heatid="20002" number="2" />
                <HEAT daytime="11:46" heatid="30002" number="3" />
                <HEAT daytime="11:48" heatid="40002" number="4" />
                <HEAT daytime="11:51" heatid="50002" number="5" />
                <HEAT daytime="11:53" heatid="60002" number="6" />
              </HEATS>
            </EVENT>
            <EVENT eventid="3" number="3" preveventid="-1" gender="M" round="PRE" daytime="11:44">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="11:57" heatid="10003" number="1" />
                <HEAT daytime="12:00" heatid="20003" number="2" />
                <HEAT daytime="12:03" heatid="30003" number="3" />
                <HEAT daytime="12:05" heatid="40003" number="4" />
                <HEAT daytime="12:07" heatid="50003" number="5" />
                <HEAT daytime="12:10" heatid="60003" number="6" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4" number="4" preveventid="-1" gender="F" round="PRE" daytime="11:59">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="12:13" heatid="10004" number="1" />
                <HEAT daytime="12:14" heatid="20004" number="2" />
                <HEAT daytime="12:17" heatid="30004" number="3" />
                <HEAT daytime="12:18" heatid="40004" number="4" />
                <HEAT daytime="12:20" heatid="50004" number="5" />
                <HEAT daytime="12:22" heatid="60004" number="6" />
              </HEATS>
            </EVENT>
            <EVENT eventid="5" number="5" preveventid="-1" gender="M" round="PRE" daytime="12:12">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="12:24" heatid="10005" number="1" />
                <HEAT daytime="12:26" heatid="20005" number="2" />
                <HEAT daytime="12:28" heatid="30005" number="3" />
                <HEAT daytime="12:30" heatid="40005" number="4" />
                <HEAT daytime="12:32" heatid="50005" number="5" />
                <HEAT daytime="12:34" heatid="60005" number="6" />
                <HEAT daytime="12:35" heatid="70005" number="7" />
                <HEAT daytime="12:37" heatid="80005" number="8" />
                <HEAT daytime="12:39" heatid="90005" number="9" />
                <HEAT daytime="12:41" heatid="100005" number="10" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6" number="6" preveventid="-1" gender="F" round="PRE" daytime="12:32">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="12:44" heatid="10006" number="1" />
                <HEAT daytime="12:48" heatid="20006" number="2" />
                <HEAT daytime="12:51" heatid="30006" number="3" />
                <HEAT daytime="12:55" heatid="40006" number="4" />
                <HEAT daytime="12:58" heatid="50006" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="7" number="7" preveventid="-1" gender="M" round="PRE" daytime="12:51">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="13:03" heatid="10007" number="1" />
                <HEAT daytime="13:06" heatid="20007" number="2" />
                <HEAT daytime="13:10" heatid="30007" number="3" />
                <HEAT daytime="13:13" heatid="40007" number="4" />
                <HEAT daytime="13:16" heatid="50007" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="8" number="8" preveventid="-1" gender="F" round="PRE" daytime="13:09">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:21" heatid="10008" number="1" />
                <HEAT daytime="13:27" heatid="20008" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9" number="9" preveventid="-1" gender="M" round="PRE" daytime="13:20">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:34" heatid="10009" number="1" />
                <HEAT daytime="13:40" heatid="20009" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="304" number="4" preveventid="4" gender="F" round="SOP" daytime="13:31">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="13:45" heatid="10304" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="305" number="5" preveventid="5" gender="M" round="SOP" daytime="13:33">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="13:47" heatid="10305" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10" number="10" preveventid="-1" gender="M" round="TIM" daytime="13:36">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:49" heatid="10010" number="1" />
                <HEAT daytime="14:07" heatid="20010" number="2" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="2" date="2022-12-13" daytime="19:30">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="101" number="1" preveventid="1" gender="F" round="FIN" daytime="19:35">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="19:38" heatid="10101" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="204" number="4" preveventid="4" gender="F" round="SEM" daytime="19:45">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="19:48" heatid="10204" number="1" />
                <HEAT daytime="19:53" heatid="20204" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="205" number="5" preveventid="5" gender="M" round="SEM" daytime="19:55">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="19:59" heatid="10205" number="1" />
                <HEAT daytime="20:03" heatid="20205" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="106" number="6" preveventid="6" gender="F" round="FIN" daytime="20:11">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="20:16" heatid="10106" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="107" number="7" preveventid="7" gender="M" round="FIN" daytime="20:19">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="20:23" heatid="10107" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="202" number="2" preveventid="2" gender="F" round="SEM" daytime="20:27">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:32" heatid="10202" number="1" />
                <HEAT daytime="20:37" heatid="20202" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="203" number="3" preveventid="3" gender="M" round="SEM" daytime="20:38">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:43" heatid="10203" number="1" />
                <HEAT daytime="20:49" heatid="20203" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="110" number="10" preveventid="10" gender="M" round="FHT" daytime="20:55">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:00" heatid="30110" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="108" number="8" preveventid="8" gender="F" round="FIN" daytime="21:22">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:25" heatid="10108" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="109" number="9" preveventid="9" gender="M" round="FIN" daytime="21:32">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:35" heatid="10109" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="3" date="2022-12-14" daytime="11:05">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="405" number="5" preveventid="205" gender="M" round="SOS" daytime="10:55">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="10:52" heatid="10405" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="11" number="11" preveventid="-1" gender="X" round="PRE" daytime="11:05">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="11:06" heatid="10011" number="1" />
                <HEAT daytime="11:10" heatid="20011" number="2" />
                <HEAT daytime="11:15" heatid="30011" number="3" />
                <HEAT daytime="11:19" heatid="40011" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="12" number="12" preveventid="-1" gender="F" round="TIM" daytime="11:19">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="11:24" heatid="10012" number="1" />
                <HEAT daytime="11:34" heatid="20012" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="13" number="13" preveventid="-1" gender="F" round="PRE" daytime="11:41">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="11:45" heatid="10013" number="1" />
                <HEAT daytime="11:48" heatid="20013" number="2" />
                <HEAT daytime="11:50" heatid="30013" number="3" />
                <HEAT daytime="11:52" heatid="40013" number="4" />
                <HEAT daytime="11:54" heatid="50013" number="5" />
                <HEAT daytime="11:56" heatid="60013" number="6" />
                <HEAT daytime="11:59" heatid="70013" number="7" />
                <HEAT daytime="12:01" heatid="80013" number="8" />
                <HEAT daytime="12:03" heatid="90013" number="9" />
              </HEATS>
            </EVENT>
            <EVENT eventid="14" number="14" preveventid="-1" gender="M" round="PRE" daytime="12:03">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:07" heatid="10014" number="1" />
                <HEAT daytime="12:10" heatid="20014" number="2" />
                <HEAT daytime="12:12" heatid="30014" number="3" />
                <HEAT daytime="12:14" heatid="40014" number="4" />
                <HEAT daytime="12:16" heatid="50014" number="5" />
                <HEAT daytime="12:18" heatid="60014" number="6" />
                <HEAT daytime="12:20" heatid="70014" number="7" />
                <HEAT daytime="12:22" heatid="80014" number="8" />
                <HEAT daytime="12:24" heatid="90014" number="9" />
                <HEAT daytime="12:26" heatid="100014" number="10" />
                <HEAT daytime="12:28" heatid="110014" number="11" />
              </HEATS>
            </EVENT>
            <EVENT eventid="15" number="15" preveventid="-1" gender="F" round="PRE" daytime="12:30">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="12:34" heatid="10015" number="1" />
                <HEAT daytime="12:37" heatid="20015" number="2" />
                <HEAT daytime="12:39" heatid="30015" number="3" />
                <HEAT daytime="12:42" heatid="40015" number="4" />
                <HEAT daytime="12:44" heatid="50015" number="5" />
                <HEAT daytime="12:47" heatid="60015" number="6" />
                <HEAT daytime="12:49" heatid="70015" number="7" />
              </HEATS>
            </EVENT>
            <EVENT eventid="16" number="16" preveventid="-1" gender="M" round="PRE" daytime="12:50">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="12:53" heatid="10016" number="1" />
                <HEAT daytime="12:55" heatid="20016" number="2" />
                <HEAT daytime="12:58" heatid="30016" number="3" />
                <HEAT daytime="13:00" heatid="40016" number="4" />
                <HEAT daytime="13:03" heatid="50016" number="5" />
                <HEAT daytime="13:05" heatid="60016" number="6" />
                <HEAT daytime="13:07" heatid="70016" number="7" />
                <HEAT daytime="13:10" heatid="80016" number="8" />
              </HEATS>
            </EVENT>
            <EVENT eventid="17" number="17" preveventid="-1" gender="F" round="PRE" daytime="13:10">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:14" heatid="10017" number="1" />
                <HEAT daytime="13:24" heatid="20017" number="2" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="4" date="2022-12-14" daytime="19:30">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="111" number="11" preveventid="11" gender="X" round="FIN" daytime="19:35">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="19:38" heatid="10111" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="112" number="12" preveventid="12" gender="F" round="FHT" daytime="19:42">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="19:47" heatid="30112" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="213" number="13" preveventid="13" gender="F" round="SEM" daytime="19:57">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="20:01" heatid="10213" number="1" />
                <HEAT daytime="20:05" heatid="20213" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="214" number="14" preveventid="14" gender="M" round="SEM" daytime="20:08">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="20:10" heatid="10214" number="1" />
                <HEAT daytime="20:16" heatid="20214" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="102" number="2" preveventid="202" gender="F" round="FIN" daytime="20:25">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:29" heatid="10102" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="103" number="3" preveventid="203" gender="M" round="FIN" daytime="20:32">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:36" heatid="10103" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="215" number="15" preveventid="15" gender="F" round="SEM" daytime="20:45">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="20:48" heatid="10215" number="1" />
                <HEAT daytime="20:54" heatid="20215" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="216" number="16" preveventid="16" gender="M" round="SEM" daytime="20:57">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="21:00" heatid="10216" number="1" />
                <HEAT daytime="21:05" heatid="20216" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="104" number="4" preveventid="204" gender="F" round="FIN" daytime="21:14">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="21:17" heatid="10104" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="105" number="5" preveventid="205" gender="M" round="FIN" daytime="21:20">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="21:23" heatid="10105" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="117" number="17" preveventid="17" gender="F" round="FIN" daytime="21:32">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:36" heatid="10117" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="5" date="2022-12-15" daytime="11:05">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="18" number="18" preveventid="-1" gender="F" round="PRE" daytime="11:05">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="11:06" heatid="10018" number="1" />
                <HEAT daytime="11:08" heatid="20018" number="2" />
                <HEAT daytime="11:10" heatid="30018" number="3" />
                <HEAT daytime="11:11" heatid="40018" number="4" />
                <HEAT daytime="11:13" heatid="50018" number="5" />
                <HEAT daytime="11:15" heatid="60018" number="6" />
                <HEAT daytime="11:17" heatid="70018" number="7" />
              </HEATS>
            </EVENT>
            <EVENT eventid="19" number="19" preveventid="-1" gender="M" round="PRE" daytime="11:19">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="11:21" heatid="10019" number="1" />
                <HEAT daytime="11:22" heatid="20019" number="2" />
                <HEAT daytime="11:25" heatid="30019" number="3" />
                <HEAT daytime="11:28" heatid="40019" number="4" />
                <HEAT daytime="11:30" heatid="50019" number="5" />
                <HEAT daytime="11:32" heatid="60019" number="6" />
              </HEATS>
            </EVENT>
            <EVENT eventid="20" number="20" preveventid="-1" gender="F" round="PRE" daytime="11:31">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="11:35" heatid="10020" number="1" />
                <HEAT daytime="11:39" heatid="20020" number="2" />
                <HEAT daytime="11:43" heatid="30020" number="3" />
                <HEAT daytime="11:46" heatid="40020" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="21" number="21" preveventid="-1" gender="M" round="PRE" daytime="11:46">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="11:50" heatid="10021" number="1" />
                <HEAT daytime="11:54" heatid="20021" number="2" />
                <HEAT daytime="11:57" heatid="30021" number="3" />
                <HEAT daytime="12:01" heatid="40021" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="22" number="22" preveventid="-1" gender="F" round="PRE" daytime="12:02">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="12:05" heatid="10022" number="1" />
                <HEAT daytime="12:07" heatid="20022" number="2" />
                <HEAT daytime="12:09" heatid="30022" number="3" />
                <HEAT daytime="12:12" heatid="40022" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="23" number="23" preveventid="-1" gender="M" round="PRE" daytime="12:12">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="12:15" heatid="10023" number="1" />
                <HEAT daytime="12:18" heatid="20023" number="2" />
                <HEAT daytime="12:20" heatid="30023" number="3" />
                <HEAT daytime="12:22" heatid="40023" number="4" />
                <HEAT daytime="12:25" heatid="50023" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="24" number="24" preveventid="-1" gender="M" round="PRE" daytime="12:25">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:28" heatid="10024" number="1" />
                <HEAT daytime="12:34" heatid="20024" number="2" />
                <HEAT daytime="12:40" heatid="30024" number="3" />
                <HEAT daytime="12:45" heatid="40024" number="4" />
                <HEAT daytime="12:50" heatid="50024" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="25" number="25" preveventid="-1" gender="F" round="PRE" daytime="12:52">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:56" heatid="10025" number="1" />
                <HEAT daytime="13:00" heatid="20025" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="26" number="26" preveventid="-1" gender="M" round="PRE" daytime="12:59">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:04" heatid="10026" number="1" />
                <HEAT daytime="13:08" heatid="20026" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="323" number="23" preveventid="23" gender="M" round="SOP" daytime="13:13">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="13:13" heatid="10323" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="6" date="2022-12-15" daytime="19:30">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="113" number="13" preveventid="213" gender="F" round="FIN" daytime="19:35">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="19:38" heatid="10113" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="114" number="14" preveventid="214" gender="M" round="FIN" daytime="19:42">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="19:45" heatid="10114" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="218" number="18" preveventid="18" gender="F" round="SEM" daytime="19:48">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="19:52" heatid="10218" number="1" />
                <HEAT daytime="19:57" heatid="20218" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="219" number="19" preveventid="19" gender="M" round="SEM" daytime="19:59">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:02" heatid="10219" number="1" />
                <HEAT daytime="20:07" heatid="20219" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="120" number="20" preveventid="20" gender="F" round="FIN" daytime="20:14">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="20:19" heatid="10120" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="121" number="21" preveventid="21" gender="M" round="FIN" daytime="20:23">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="20:28" heatid="10121" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="115" number="15" preveventid="215" gender="F" round="FIN" daytime="20:37">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="20:42" heatid="10115" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="116" number="16" preveventid="216" gender="M" round="FIN" daytime="20:44">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="20:49" heatid="10116" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="222" number="22" preveventid="22" gender="F" round="SEM" daytime="20:57">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="21:00" heatid="10222" number="1" />
                <HEAT daytime="21:06" heatid="20222" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="223" number="23" preveventid="23" gender="M" round="SEM" daytime="21:14">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="21:17" heatid="10223" number="1" />
                <HEAT daytime="21:23" heatid="20223" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="124" number="24" preveventid="24" gender="M" round="FIN" daytime="21:31">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:35" heatid="10124" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="125" number="25" preveventid="25" gender="F" round="FIN" daytime="21:46">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:51" heatid="10125" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="126" number="26" preveventid="26" gender="M" round="FIN" daytime="21:54">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:58" heatid="10126" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="7" date="2022-12-16" daytime="11:05">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="27" number="27" preveventid="-1" gender="X" round="PRE" daytime="11:05">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="11:06" heatid="10027" number="1" />
                <HEAT daytime="11:10" heatid="20027" number="2" />
                <HEAT daytime="11:14" heatid="30027" number="3" />
                <HEAT daytime="11:17" heatid="40027" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="28" number="28" preveventid="-1" gender="F" round="PRE" daytime="11:19">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="11:21" heatid="10028" number="1" />
                <HEAT daytime="11:25" heatid="20028" number="2" />
                <HEAT daytime="11:28" heatid="30028" number="3" />
                <HEAT daytime="11:32" heatid="40028" number="4" />
                <HEAT daytime="11:36" heatid="50028" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="29" number="29" preveventid="-1" gender="M" round="PRE" daytime="11:39">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="11:41" heatid="10029" number="1" />
                <HEAT daytime="11:45" heatid="20029" number="2" />
                <HEAT daytime="11:49" heatid="30029" number="3" />
                <HEAT daytime="11:53" heatid="40029" number="4" />
                <HEAT daytime="11:56" heatid="50029" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="30" number="30" preveventid="-1" gender="F" round="PRE" daytime="11:58">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:00" heatid="10030" number="1" />
                <HEAT daytime="12:02" heatid="20030" number="2" />
                <HEAT daytime="12:04" heatid="30030" number="3" />
                <HEAT daytime="12:05" heatid="40030" number="4" />
                <HEAT daytime="12:07" heatid="50030" number="5" />
                <HEAT daytime="12:09" heatid="60030" number="6" />
                <HEAT daytime="12:10" heatid="70030" number="7" />
                <HEAT daytime="12:12" heatid="80030" number="8" />
              </HEATS>
            </EVENT>
            <EVENT eventid="31" number="31" preveventid="-1" gender="M" round="PRE" daytime="12:14">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:16" heatid="10031" number="1" />
                <HEAT daytime="12:17" heatid="20031" number="2" />
                <HEAT daytime="12:19" heatid="30031" number="3" />
                <HEAT daytime="12:20" heatid="40031" number="4" />
                <HEAT daytime="12:22" heatid="50031" number="5" />
                <HEAT daytime="12:24" heatid="60031" number="6" />
                <HEAT daytime="12:26" heatid="70031" number="7" />
                <HEAT daytime="12:27" heatid="80031" number="8" />
                <HEAT daytime="12:29" heatid="90031" number="9" />
                <HEAT daytime="12:31" heatid="100031" number="10" />
                <HEAT daytime="12:33" heatid="110031" number="11" />
              </HEATS>
            </EVENT>
            <EVENT eventid="32" number="32" preveventid="-1" gender="M" round="PRE" daytime="12:36">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:36" heatid="10032" number="1" />
                <HEAT daytime="12:45" heatid="20032" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="419" number="19" preveventid="219" gender="M" round="SOS" daytime="12:55">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="12:55" heatid="10419" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="33" number="33" preveventid="-1" gender="F" round="TIM" daytime="12:57">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="12:58" heatid="10033" number="1" />
                <HEAT daytime="13:16" heatid="20033" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="331" number="31" preveventid="31" gender="M" round="SOP" daytime="13:35">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:36" heatid="10331" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="8" date="2022-12-16" daytime="19:30">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="127" number="27" preveventid="27" gender="X" round="FIN" daytime="19:35">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="19:38" heatid="10127" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="128" number="28" preveventid="28" gender="F" round="FIN" daytime="19:42">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="19:45" heatid="10128" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="129" number="29" preveventid="29" gender="M" round="FIN" daytime="19:51">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="19:54" heatid="10129" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="118" number="18" preveventid="218" gender="F" round="FIN" daytime="20:06">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:10" heatid="10118" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="230" number="30" preveventid="30" gender="F" round="SEM" daytime="20:25">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="20:29" heatid="10230" number="1" />
                <HEAT daytime="20:33" heatid="20230" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="231" number="31" preveventid="31" gender="M" round="SEM" daytime="20:41">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="20:44" heatid="10231" number="1" />
                <HEAT daytime="20:49" heatid="20231" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="122" number="22" preveventid="222" gender="F" round="FIN" daytime="20:56">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="20:59" heatid="10122" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="123" number="23" preveventid="223" gender="M" round="FIN" daytime="21:04">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="21:06" heatid="10123" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="119" number="19" preveventid="219" gender="M" round="FIN" daytime="21:11">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="21:14" heatid="10119" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="133" number="33" preveventid="33" gender="F" round="FHT" daytime="21:16">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:20" heatid="30133" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="132" number="32" preveventid="32" gender="M" round="FIN" daytime="21:45">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:49" heatid="10132" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="9" date="2022-12-17" daytime="11:05">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="34" number="34" preveventid="-1" gender="F" round="PRE" daytime="11:05">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="11:06" heatid="10034" number="1" />
                <HEAT daytime="11:10" heatid="20034" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="35" number="35" preveventid="-1" gender="M" round="PRE" daytime="11:12">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="11:15" heatid="10035" number="1" />
                <HEAT daytime="11:19" heatid="20035" number="2" />
                <HEAT daytime="11:23" heatid="30035" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="36" number="36" preveventid="-1" gender="F" round="PRE" daytime="11:21">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="11:27" heatid="10036" number="1" />
                <HEAT daytime="11:33" heatid="20036" number="2" />
                <HEAT daytime="11:39" heatid="30036" number="3" />
                <HEAT daytime="11:45" heatid="40036" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="37" number="37" preveventid="-1" gender="M" round="PRE" daytime="11:47">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="11:52" heatid="10037" number="1" />
                <HEAT daytime="11:58" heatid="20037" number="2" />
                <HEAT daytime="12:04" heatid="30037" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="38" number="38" preveventid="-1" gender="F" round="PRE" daytime="12:05">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="12:10" heatid="10038" number="1" />
                <HEAT daytime="12:12" heatid="20038" number="2" />
                <HEAT daytime="12:15" heatid="30038" number="3" />
                <HEAT daytime="12:17" heatid="40038" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="39" number="39" preveventid="-1" gender="M" round="PRE" daytime="12:16">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="12:20" heatid="10039" number="1" />
                <HEAT daytime="12:22" heatid="20039" number="2" />
                <HEAT daytime="12:25" heatid="30039" number="3" />
                <HEAT daytime="12:27" heatid="40039" number="4" />
                <HEAT daytime="12:29" heatid="50039" number="5" />
                <HEAT daytime="12:34" heatid="60039" number="6" />
                <HEAT daytime="12:37" heatid="70039" number="7" />
                <HEAT daytime="12:39" heatid="80039" number="8" />
              </HEATS>
            </EVENT>
            <EVENT eventid="40" number="40" preveventid="-1" gender="F" round="PRE" daytime="12:36">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="12:43" heatid="10040" number="1" />
                <HEAT daytime="12:45" heatid="20040" number="2" />
                <HEAT daytime="12:47" heatid="30040" number="3" />
                <HEAT daytime="12:48" heatid="40040" number="4" />
                <HEAT daytime="12:51" heatid="50040" number="5" />
                <HEAT daytime="12:53" heatid="60040" number="6" />
                <HEAT daytime="12:55" heatid="70040" number="7" />
              </HEATS>
            </EVENT>
            <EVENT eventid="41" number="41" preveventid="-1" gender="M" round="PRE" daytime="12:51">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="12:58" heatid="10041" number="1" />
                <HEAT daytime="13:00" heatid="20041" number="2" />
                <HEAT daytime="13:01" heatid="30041" number="3" />
                <HEAT daytime="13:04" heatid="40041" number="4" />
                <HEAT daytime="13:05" heatid="50041" number="5" />
                <HEAT daytime="13:08" heatid="60041" number="6" />
                <HEAT daytime="13:11" heatid="70041" number="7" />
                <HEAT daytime="13:13" heatid="80041" number="8" />
                <HEAT daytime="13:16" heatid="90041" number="9" />
              </HEATS>
            </EVENT>
            <EVENT eventid="338" number="38" preveventid="38" gender="F" round="SOP" daytime="13:09">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="13:20" heatid="10338" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="42" number="42" preveventid="-1" gender="M" round="TIM" daytime="13:12">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="13:22" heatid="10042" number="1" />
                <HEAT daytime="13:32" heatid="20042" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="341" number="41" preveventid="41" gender="M" round="SOP" daytime="13:33">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="13:42" heatid="10341" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="10" date="2022-12-17" daytime="19:30">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="134" number="34" preveventid="34" gender="F" round="FIN" daytime="19:35">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="19:38" heatid="10134" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="135" number="35" preveventid="35" gender="M" round="FIN" daytime="19:43">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="19:46" heatid="10135" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="142" number="42" preveventid="42" gender="M" round="FHT" daytime="19:50">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="19:55" heatid="30142" number="3" />
              </HEATS>
            </EVENT>
            <EVENT eventid="238" number="38" preveventid="38" gender="F" round="SEM" daytime="20:11">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="20:15" heatid="10238" number="1" />
                <HEAT daytime="20:20" heatid="20238" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="239" number="39" preveventid="39" gender="M" round="SEM" daytime="20:22">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="20:26" heatid="10239" number="1" />
                <HEAT daytime="20:31" heatid="20239" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="136" number="36" preveventid="36" gender="F" round="FIN" daytime="20:40">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="20:45" heatid="10136" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="137" number="37" preveventid="37" gender="M" round="FIN" daytime="20:50">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="20:56" heatid="10137" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="240" number="40" preveventid="40" gender="F" round="SEM" daytime="21:07">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="21:11" heatid="10240" number="1" />
                <HEAT daytime="21:15" heatid="20240" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="241" number="41" preveventid="41" gender="M" round="SEM" daytime="21:17">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="21:22" heatid="10241" number="1" />
                <HEAT daytime="21:26" heatid="20241" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="130" number="30" preveventid="230" gender="F" round="FIN" daytime="21:33">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:37" heatid="10130" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="131" number="31" preveventid="231" gender="M" round="FIN" daytime="21:39">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="21:43" heatid="10131" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="11" date="2022-12-18" daytime="11:05">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="43" number="43" preveventid="-1" gender="F" round="PRE" daytime="11:05">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="11:06" heatid="10043" number="1" />
                <HEAT daytime="11:09" heatid="20043" number="2" />
                <HEAT daytime="11:13" heatid="30043" number="3" />
                <HEAT daytime="11:16" heatid="40043" number="4" />
                <HEAT daytime="11:20" heatid="50043" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="44" number="44" preveventid="-1" gender="M" round="PRE" daytime="11:23">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="11:24" heatid="10044" number="1" />
                <HEAT daytime="11:27" heatid="20044" number="2" />
                <HEAT daytime="11:30" heatid="30044" number="3" />
                <HEAT daytime="11:33" heatid="40044" number="4" />
                <HEAT daytime="11:36" heatid="50044" number="5" />
                <HEAT daytime="11:40" heatid="60044" number="6" />
              </HEATS>
            </EVENT>
            <EVENT eventid="45" number="45" preveventid="-1" gender="F" round="PRE" daytime="11:44">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="11:44" heatid="10045" number="1" />
                <HEAT daytime="11:48" heatid="20045" number="2" />
                <HEAT daytime="11:52" heatid="30045" number="3" />
                <HEAT daytime="11:55" heatid="40045" number="4" />
                <HEAT daytime="11:59" heatid="50045" number="5" />
              </HEATS>
            </EVENT>
            <EVENT eventid="46" number="46" preveventid="-1" gender="M" round="PRE" daytime="12:03">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="12:03" heatid="10046" number="1" />
                <HEAT daytime="12:07" heatid="20046" number="2" />
                <HEAT daytime="12:10" heatid="30046" number="3" />
                <HEAT daytime="12:14" heatid="40046" number="4" />
              </HEATS>
            </EVENT>
            <EVENT eventid="47" number="47" preveventid="-1" gender="F" round="PRE" daytime="12:17">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="12:18" heatid="10047" number="1" />
                <HEAT daytime="12:25" heatid="20047" number="2" />
              </HEATS>
            </EVENT>
            <EVENT eventid="48" number="48" preveventid="-1" gender="M" round="PRE" daytime="12:29">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="12:32" heatid="10048" number="1" />
                <HEAT daytime="12:38" heatid="20048" number="2" />
                <HEAT daytime="12:44" heatid="30048" number="3" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION number="12" date="2022-12-18" daytime="19:30">
          <POOL lanemax="9" lanemin="1" />
          <EVENTS>
            <EVENT eventid="138" number="38" preveventid="238" gender="F" round="FIN" daytime="19:35">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="19:38" heatid="10138" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="139" number="39" preveventid="239" gender="M" round="FIN" daytime="19:42">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <HEATS>
                <HEAT daytime="19:45" heatid="10139" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="140" number="40" preveventid="240" gender="F" round="FIN" daytime="19:49">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="19:52" heatid="10140" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="141" number="41" preveventid="241" gender="M" round="FIN" daytime="20:01">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT daytime="20:04" heatid="10141" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="145" number="45" preveventid="45" gender="F" round="FIN" daytime="20:08">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:11" heatid="10145" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="146" number="46" preveventid="46" gender="M" round="FIN" daytime="20:22">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <HEATS>
                <HEAT daytime="20:26" heatid="10146" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="143" number="43" preveventid="43" gender="F" round="FIN" daytime="20:36">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="20:39" heatid="10143" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="144" number="44" preveventid="44" gender="M" round="FIN" daytime="20:50">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT daytime="20:53" heatid="10144" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="147" number="47" preveventid="47" gender="F" round="FIN" daytime="21:03">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="21:09" heatid="10147" number="1" />
              </HEATS>
            </EVENT>
            <EVENT eventid="148" number="48" preveventid="48" gender="M" round="FIN" daytime="21:19">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <HEATS>
                <HEAT daytime="21:27" heatid="10148" number="1" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB name="Afghanistan" shortname="AFG" code="AFG" nation="AFG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="164222" lastname="ANWARI" firstname="Fahim" gender="M" birthdate="1999-05-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.52" eventid="5" heat="3" lane="1">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.67" eventid="31" heat="3" lane="8">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="62" lane="1" heat="3" heatid="30005" swimtime="00:00:28.48" reactiontime="+67" points="445">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.23" />
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="74" lane="8" heat="3" heatid="30031" swimtime="00:00:27.30" reactiontime="+74" points="402">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Albania" shortname="ALB" code="ALB" nation="ALB" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="162857" lastname="PRISKA" firstname="Paolo" gender="M" birthdate="2004-09-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.05" eventid="39" heat="2" lane="5">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.14" eventid="14" heat="4" lane="7">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="49" lane="5" heat="2" heatid="20039" swimtime="00:00:57.30" reactiontime="+60" points="579">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:26.89" />
                    <SPLIT distance="75" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:00:57.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="64" lane="7" heat="4" heatid="40014" swimtime="00:00:52.18" reactiontime="+63" points="634">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:24.89" />
                    <SPLIT distance="75" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213756" lastname="DUCAJ" firstname="Mark" gender="M" birthdate="2003-05-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.08" eventid="44" heat="2" lane="7">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:03:58.97" eventid="24" heat="1" lane="3">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="38" lane="7" heat="2" heatid="20044" swimtime="00:01:50.38" reactiontime="+71" points="729">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:25.74" />
                    <SPLIT distance="75" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:00:53.72" />
                    <SPLIT distance="125" swimtime="00:01:07.89" />
                    <SPLIT distance="150" swimtime="00:01:21.97" />
                    <SPLIT distance="175" swimtime="00:01:36.43" />
                    <SPLIT distance="200" swimtime="00:01:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="29" lane="3" heat="1" heatid="10024" swimtime="00:03:56.41" reactiontime="+78" points="723">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="75" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:00:55.99" />
                    <SPLIT distance="125" swimtime="00:01:11.01" />
                    <SPLIT distance="150" swimtime="00:01:25.91" />
                    <SPLIT distance="175" swimtime="00:01:40.92" />
                    <SPLIT distance="200" swimtime="00:01:55.89" />
                    <SPLIT distance="225" swimtime="00:02:11.12" />
                    <SPLIT distance="250" swimtime="00:02:26.36" />
                    <SPLIT distance="275" swimtime="00:02:41.52" />
                    <SPLIT distance="300" swimtime="00:02:56.79" />
                    <SPLIT distance="325" swimtime="00:03:12.12" />
                    <SPLIT distance="350" swimtime="00:03:27.31" />
                    <SPLIT distance="375" swimtime="00:03:42.33" />
                    <SPLIT distance="400" swimtime="00:03:56.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213888" lastname="MECA" firstname="Kaltra" gender="F" birthdate="2008-03-26">
              <ENTRIES>
                <ENTRY entrytime="00:02:15.56" eventid="43" heat="1" lane="3">
                  <MEETINFO date="2022-07-26" />
                </ENTRY>
                <ENTRY entrytime="00:04:37.39" eventid="1" heat="1" lane="2">
                  <MEETINFO date="2022-07-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="31" lane="3" heat="1" heatid="10043" swimtime="00:02:10.75" reactiontime="+81" points="600">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.60" />
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="75" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:03.03" />
                    <SPLIT distance="125" swimtime="00:01:19.90" />
                    <SPLIT distance="150" swimtime="00:01:37.11" />
                    <SPLIT distance="175" swimtime="00:01:54.22" />
                    <SPLIT distance="200" swimtime="00:02:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="27" lane="2" heat="1" heatid="10001" swimtime="00:04:31.99" reactiontime="+90" points="636">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="75" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:02.60" />
                    <SPLIT distance="125" swimtime="00:01:19.52" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                    <SPLIT distance="175" swimtime="00:01:54.29" />
                    <SPLIT distance="200" swimtime="00:02:11.59" />
                    <SPLIT distance="225" swimtime="00:02:29.06" />
                    <SPLIT distance="250" swimtime="00:02:46.61" />
                    <SPLIT distance="275" swimtime="00:03:04.07" />
                    <SPLIT distance="300" swimtime="00:03:21.80" />
                    <SPLIT distance="325" swimtime="00:03:39.54" />
                    <SPLIT distance="350" swimtime="00:03:57.46" />
                    <SPLIT distance="375" swimtime="00:04:15.10" />
                    <SPLIT distance="400" swimtime="00:04:31.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Algeria" shortname="ALG" code="ALG" nation="ALG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="149785" lastname="ARDJOUNE" firstname="Abdellah" gender="M" birthdate="2001-02-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.31" eventid="3" heat="2" lane="5">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.88" eventid="46" heat="1" lane="4">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.78" eventid="19" heat="1" lane="4">
                  <MEETINFO date="2021-10-11" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="36" lane="5" heat="2" heatid="20003" swimtime="00:00:55.54" reactiontime="+67" points="658">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:00:55.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="23" lane="4" heat="1" heatid="10046" swimtime="00:01:59.78" reactiontime="+62" points="685">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="75" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:00:57.47" />
                    <SPLIT distance="125" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:28.76" />
                    <SPLIT distance="175" swimtime="00:01:44.55" />
                    <SPLIT distance="200" swimtime="00:01:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="36" lane="4" heat="1" heatid="10019" swimtime="00:00:25.71" reactiontime="+66" points="645">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113400" lastname="MELIH" firstname="Amel" gender="F" birthdate="1993-10-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.34" eventid="13" heat="5" lane="4">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.77" eventid="30" heat="4" lane="4">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="36" lane="4" heat="5" heatid="50013" swimtime="00:00:55.58" reactiontime="+62" points="739">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.46" />
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="75" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:00:55.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="26" lane="4" heat="4" heatid="40030" swimtime="00:00:25.09" reactiontime="+60" points="763">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.27" />
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Andorra" shortname="AND" code="AND" nation="AND" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154153" lastname="LOMERO ARENAS" firstname="Tomàs" gender="M" birthdate="2001-07-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.48" eventid="39" heat="3" lane="2">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:50.42" eventid="14" heat="5" lane="3">
                  <MEETINFO date="2021-11-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="40" lane="2" heat="3" heatid="30039" swimtime="00:00:54.01" reactiontime="+60" points="692">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.33" />
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="75" swimtime="00:00:38.99" />
                    <SPLIT distance="100" swimtime="00:00:54.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="53" lane="3" heat="5" heatid="50014" swimtime="00:00:50.32" reactiontime="+61" points="707">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:23.95" />
                    <SPLIT distance="75" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:00:50.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128785" lastname="LOMERO" firstname="Bernat" gender="M" birthdate="1997-12-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.33" eventid="5" heat="4" lane="6">
                  <MEETINFO date="2022-04-13" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.67" eventid="31" heat="6" lane="8">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="51" lane="6" heat="4" heatid="40005" swimtime="00:00:24.29" reactiontime="+63" points="717">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.88" />
                    <SPLIT distance="50" swimtime="00:00:24.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="51" lane="8" heat="6" heatid="60031" swimtime="00:00:22.93" reactiontime="+62" points="679">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.97" />
                    <SPLIT distance="50" swimtime="00:00:22.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105101" lastname="TUDO CUBELLS" firstname="Nadia" gender="F" birthdate="1997-04-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:10.70" eventid="15" heat="3" lane="2">
                  <MEETINFO date="2021-10-02" />
                </ENTRY>
                <ENTRY entrytime="00:02:30.40" eventid="28" heat="1" lane="4">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="39" lane="2" heat="3" heatid="30015" swimtime="00:01:11.31" reactiontime="+68" points="668">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.57" />
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="75" swimtime="00:00:52.34" />
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="28" lane="4" heat="1" heatid="10028" swimtime="00:02:31.45" reactiontime="+67" points="701">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.79" />
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="75" swimtime="00:00:53.22" />
                    <SPLIT distance="100" swimtime="00:01:12.67" />
                    <SPLIT distance="125" swimtime="00:01:32.35" />
                    <SPLIT distance="150" swimtime="00:01:52.01" />
                    <SPLIT distance="175" swimtime="00:02:11.66" />
                    <SPLIT distance="200" swimtime="00:02:31.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Antigua &amp; Barbuda" shortname="ANT" code="ANT" nation="ANT" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="150205" lastname="WUILLIEZ" firstname="Jadon" gender="M" birthdate="2002-06-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.73" eventid="16" heat="5" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.98" eventid="41" heat="6" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="39" lane="8" heat="5" heatid="50016" swimtime="00:01:00.00" reactiontime="+67" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.46" />
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="75" swimtime="00:00:43.63" />
                    <SPLIT distance="100" swimtime="00:01:00.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="30" lane="2" heat="6" heatid="60041" swimtime="00:00:27.16" reactiontime="+64" points="775">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Argentina" shortname="ARG" code="ARG" nation="ARG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="147577" lastname="ALBA" firstname="Lucas Ezequiel" gender="M" birthdate="2000-09-17">
              <ENTRIES>
                <ENTRY entrytime="00:14:56.52" eventid="10" heat="2" lane="8">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:03:47.20" eventid="24" heat="3" lane="8">
                  <MEETINFO date="2022-10-20" />
                </ENTRY>
                <ENTRY entrytime="00:07:49.65" eventid="42" heat="2" lane="2">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="12" lane="8" heat="2" heatid="20010" swimtime="00:14:56.41" reactiontime="+68" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="75" swimtime="00:00:41.38" />
                    <SPLIT distance="100" swimtime="00:00:55.87" />
                    <SPLIT distance="125" swimtime="00:01:10.43" />
                    <SPLIT distance="150" swimtime="00:01:25.19" />
                    <SPLIT distance="175" swimtime="00:01:39.88" />
                    <SPLIT distance="200" swimtime="00:01:54.70" />
                    <SPLIT distance="225" swimtime="00:02:09.38" />
                    <SPLIT distance="250" swimtime="00:02:24.11" />
                    <SPLIT distance="275" swimtime="00:02:38.96" />
                    <SPLIT distance="300" swimtime="00:02:53.84" />
                    <SPLIT distance="325" swimtime="00:03:08.54" />
                    <SPLIT distance="350" swimtime="00:03:23.38" />
                    <SPLIT distance="375" swimtime="00:03:38.22" />
                    <SPLIT distance="400" swimtime="00:03:53.05" />
                    <SPLIT distance="425" swimtime="00:04:07.83" />
                    <SPLIT distance="450" swimtime="00:04:22.81" />
                    <SPLIT distance="475" swimtime="00:04:37.61" />
                    <SPLIT distance="500" swimtime="00:04:52.53" />
                    <SPLIT distance="525" swimtime="00:05:07.30" />
                    <SPLIT distance="550" swimtime="00:05:22.30" />
                    <SPLIT distance="575" swimtime="00:05:37.19" />
                    <SPLIT distance="600" swimtime="00:05:52.04" />
                    <SPLIT distance="625" swimtime="00:06:07.09" />
                    <SPLIT distance="650" swimtime="00:06:21.97" />
                    <SPLIT distance="675" swimtime="00:06:37.02" />
                    <SPLIT distance="700" swimtime="00:06:52.04" />
                    <SPLIT distance="725" swimtime="00:07:07.07" />
                    <SPLIT distance="750" swimtime="00:07:22.07" />
                    <SPLIT distance="775" swimtime="00:07:37.22" />
                    <SPLIT distance="800" swimtime="00:07:52.07" />
                    <SPLIT distance="825" swimtime="00:08:06.98" />
                    <SPLIT distance="850" swimtime="00:08:21.98" />
                    <SPLIT distance="875" swimtime="00:08:37.15" />
                    <SPLIT distance="900" swimtime="00:08:52.24" />
                    <SPLIT distance="925" swimtime="00:09:07.35" />
                    <SPLIT distance="950" swimtime="00:09:22.30" />
                    <SPLIT distance="975" swimtime="00:09:37.32" />
                    <SPLIT distance="1000" swimtime="00:09:52.23" />
                    <SPLIT distance="1025" swimtime="00:10:07.48" />
                    <SPLIT distance="1050" swimtime="00:10:22.55" />
                    <SPLIT distance="1075" swimtime="00:10:37.73" />
                    <SPLIT distance="1100" swimtime="00:10:52.80" />
                    <SPLIT distance="1125" swimtime="00:11:07.95" />
                    <SPLIT distance="1150" swimtime="00:11:23.28" />
                    <SPLIT distance="1175" swimtime="00:11:38.65" />
                    <SPLIT distance="1200" swimtime="00:11:53.80" />
                    <SPLIT distance="1225" swimtime="00:12:08.99" />
                    <SPLIT distance="1250" swimtime="00:12:24.37" />
                    <SPLIT distance="1275" swimtime="00:12:39.64" />
                    <SPLIT distance="1300" swimtime="00:12:54.89" />
                    <SPLIT distance="1325" swimtime="00:13:10.25" />
                    <SPLIT distance="1350" swimtime="00:13:25.69" />
                    <SPLIT distance="1375" swimtime="00:13:41.07" />
                    <SPLIT distance="1400" swimtime="00:13:56.37" />
                    <SPLIT distance="1425" swimtime="00:14:11.80" />
                    <SPLIT distance="1450" swimtime="00:14:27.05" />
                    <SPLIT distance="1475" swimtime="00:14:42.16" />
                    <SPLIT distance="1500" swimtime="00:14:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="23" lane="8" heat="3" heatid="30024" swimtime="00:03:48.47" reactiontime="+66" points="801">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.14" />
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="75" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:00:54.32" />
                    <SPLIT distance="125" swimtime="00:01:08.71" />
                    <SPLIT distance="150" swimtime="00:01:23.10" />
                    <SPLIT distance="175" swimtime="00:01:37.63" />
                    <SPLIT distance="200" swimtime="00:01:52.05" />
                    <SPLIT distance="225" swimtime="00:02:06.43" />
                    <SPLIT distance="250" swimtime="00:02:20.84" />
                    <SPLIT distance="275" swimtime="00:02:35.31" />
                    <SPLIT distance="300" swimtime="00:02:49.89" />
                    <SPLIT distance="325" swimtime="00:03:04.57" />
                    <SPLIT distance="350" swimtime="00:03:19.35" />
                    <SPLIT distance="375" swimtime="00:03:34.21" />
                    <SPLIT distance="400" swimtime="00:03:48.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="15" lane="2" heat="2" heatid="20042" swimtime="00:07:49.53" reactiontime="+65" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.15" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:54.56" />
                    <SPLIT distance="125" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:23.32" />
                    <SPLIT distance="175" swimtime="00:01:37.94" />
                    <SPLIT distance="200" swimtime="00:01:52.69" />
                    <SPLIT distance="225" swimtime="00:02:07.44" />
                    <SPLIT distance="250" swimtime="00:02:22.20" />
                    <SPLIT distance="275" swimtime="00:02:36.91" />
                    <SPLIT distance="300" swimtime="00:02:51.77" />
                    <SPLIT distance="325" swimtime="00:03:06.50" />
                    <SPLIT distance="350" swimtime="00:03:21.16" />
                    <SPLIT distance="375" swimtime="00:03:36.04" />
                    <SPLIT distance="400" swimtime="00:03:50.92" />
                    <SPLIT distance="425" swimtime="00:04:05.78" />
                    <SPLIT distance="450" swimtime="00:04:20.53" />
                    <SPLIT distance="475" swimtime="00:04:35.18" />
                    <SPLIT distance="500" swimtime="00:04:50.05" />
                    <SPLIT distance="525" swimtime="00:05:04.87" />
                    <SPLIT distance="550" swimtime="00:05:19.70" />
                    <SPLIT distance="575" swimtime="00:05:34.66" />
                    <SPLIT distance="600" swimtime="00:05:49.63" />
                    <SPLIT distance="625" swimtime="00:06:04.58" />
                    <SPLIT distance="650" swimtime="00:06:19.53" />
                    <SPLIT distance="675" swimtime="00:06:34.56" />
                    <SPLIT distance="700" swimtime="00:06:49.58" />
                    <SPLIT distance="725" swimtime="00:07:04.71" />
                    <SPLIT distance="750" swimtime="00:07:20.03" />
                    <SPLIT distance="775" swimtime="00:07:35.10" />
                    <SPLIT distance="800" swimtime="00:07:49.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110696" lastname="BERRINO" firstname="Andrea" gender="F" birthdate="1994-02-14">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.40" eventid="2" heat="3" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.00" eventid="45" heat="2" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.20" eventid="18" heat="6" lane="1">
                  <MEETINFO date="2022-10-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.25" eventid="30" heat="5" lane="5">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="27" lane="3" heat="3" heatid="30002" swimtime="00:00:58.85" reactiontime="+58" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="75" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:00:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="24" lane="3" heat="2" heatid="20045" swimtime="00:02:08.10" reactiontime="+57" points="800">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="75" swimtime="00:00:46.42" />
                    <SPLIT distance="100" swimtime="00:01:02.84" />
                    <SPLIT distance="125" swimtime="00:01:19.35" />
                    <SPLIT distance="150" swimtime="00:01:35.75" />
                    <SPLIT distance="175" swimtime="00:01:52.32" />
                    <SPLIT distance="200" swimtime="00:02:08.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="23" lane="1" heat="6" heatid="60018" swimtime="00:00:27.15" reactiontime="+57" points="806">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="20" lane="5" heat="5" heatid="50030" swimtime="00:00:24.93" reactiontime="+68" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125910" lastname="CEBALLOS" firstname="Macarena" gender="F" birthdate="1995-01-12">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.71" eventid="15" heat="4" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.97" eventid="28" heat="2" lane="3">
                  <MEETINFO date="2022-10-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.04" eventid="40" heat="5" lane="2">
                  <MEETINFO date="2022-09-15" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="22" lane="7" heat="4" heatid="40015" swimtime="00:01:05.62" reactiontime="+68" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.20" />
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="75" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:05.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="16" lane="3" heat="2" heatid="20028" swimtime="00:02:22.10" reactiontime="+67" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.88" />
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="75" swimtime="00:00:50.00" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="125" swimtime="00:01:26.31" />
                    <SPLIT distance="150" swimtime="00:01:44.68" />
                    <SPLIT distance="175" swimtime="00:02:03.30" />
                    <SPLIT distance="200" swimtime="00:02:22.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="16" lane="2" heat="5" heatid="50040" swimtime="00:00:30.33" reactiontime="+62" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="14" lane="8" heat="1" heatid="10240" swimtime="00:00:30.10" reactiontime="+67" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.80" />
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Armenia" shortname="ARM" code="ARM" nation="ARM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="129469" lastname="BARSEGHYAN" firstname="Artur" gender="M" birthdate="2002-03-29">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.50" eventid="5" heat="6" lane="2">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.49" eventid="31" heat="6" lane="7">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="46" lane="2" heat="6" heatid="60005" swimtime="00:00:23.65" reactiontime="+66" points="777">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.93" />
                    <SPLIT distance="50" swimtime="00:00:23.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="47" lane="7" heat="6" heatid="60031" swimtime="00:00:22.30" reactiontime="+65" points="738">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.73" />
                    <SPLIT distance="50" swimtime="00:00:22.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108147" lastname="POGHOSYAN" firstname="Ani" gender="F" birthdate="2000-06-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.58" eventid="13" heat="4" lane="6">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.14" eventid="43" heat="1" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="44" lane="6" heat="4" heatid="40013" swimtime="00:00:57.91" reactiontime="+75" points="653">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:27.53" />
                    <SPLIT distance="75" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="29" lane="4" heat="1" heatid="10043" swimtime="00:02:04.30" reactiontime="+74" points="698">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="75" swimtime="00:00:44.27" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="125" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:31.85" />
                    <SPLIT distance="175" swimtime="00:01:48.37" />
                    <SPLIT distance="200" swimtime="00:02:04.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Aruba" shortname="ARU" code="ARU" nation="ARU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="105498" lastname="SCHREUDERS" firstname="Mikel" gender="M" birthdate="1998-09-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.01" eventid="14" heat="10" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:01:46.08" eventid="44" heat="3" lane="2">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.52" eventid="41" heat="5" lane="7">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.80" eventid="31" heat="8" lane="8">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.25" eventid="23" heat="3" lane="1">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="16" lane="1" heat="10" heatid="100014" swimtime="00:00:47.03" reactiontime="+62" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.66" />
                    <SPLIT distance="50" swimtime="00:00:22.61" />
                    <SPLIT distance="75" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:00:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="15" lane="8" heat="1" heatid="10214" swimtime="00:00:47.12" reactiontime="+64" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.97" />
                    <SPLIT distance="50" swimtime="00:00:22.89" />
                    <SPLIT distance="75" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:00:47.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="35" lane="2" heat="3" heatid="30044" swimtime="00:01:47.74" reactiontime="+62" points="784">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:24.22" />
                    <SPLIT distance="75" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:00:50.89" />
                    <SPLIT distance="125" swimtime="00:01:04.69" />
                    <SPLIT distance="150" swimtime="00:01:19.03" />
                    <SPLIT distance="175" swimtime="00:01:33.57" />
                    <SPLIT distance="200" swimtime="00:01:47.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="15" lane="7" heat="5" heatid="50041" swimtime="00:00:26.47" reactiontime="+63" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="15" lane="8" heat="2" heatid="20241" swimtime="00:00:26.66" reactiontime="+64" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="38" lane="8" heat="8" heatid="80031" swimtime="00:00:21.61" reactiontime="+64" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:21.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="15" lane="1" heat="3" heatid="30023" swimtime="00:00:52.65" reactiontime="+63" points="820">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.81" />
                    <SPLIT distance="50" swimtime="00:00:24.80" />
                    <SPLIT distance="75" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:00:52.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="12" lane="8" heat="2" heatid="20223" swimtime="00:00:52.34" reactiontime="+65" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:24.67" />
                    <SPLIT distance="75" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123675" lastname="TIMMER" firstname="Elisabeth" gender="F" birthdate="2001-03-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.78" eventid="13" heat="4" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.16" eventid="30" heat="4" lane="6">
                  <MEETINFO date="2022-10-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="39" lane="7" heat="4" heatid="40013" swimtime="00:00:55.88" reactiontime="+68" points="727">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="75" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="31" lane="6" heat="4" heatid="40030" swimtime="00:00:25.64" reactiontime="+68" points="715">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.37" />
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Australia" shortname="AUS" code="AUS" nation="AUS" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="120897" lastname="WOODWARD" firstname="Bradley" gender="M" birthdate="1998-07-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.10" eventid="3" heat="6" lane="7">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.14" eventid="46" heat="2" lane="6">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.08" eventid="19" heat="3" lane="1">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="22" lane="7" heat="6" heatid="60003" swimtime="00:00:51.35" reactiontime="+66" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:24.87" />
                    <SPLIT distance="75" swimtime="00:00:38.21" />
                    <SPLIT distance="100" swimtime="00:00:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="9" lane="6" heat="2" heatid="20046" swimtime="00:01:51.46" reactiontime="+64" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                    <SPLIT distance="50" swimtime="00:00:26.18" />
                    <SPLIT distance="75" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:00:54.41" />
                    <SPLIT distance="125" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:22.86" />
                    <SPLIT distance="175" swimtime="00:01:37.44" />
                    <SPLIT distance="200" swimtime="00:01:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="23" lane="1" heat="3" heatid="30019" swimtime="00:00:23.80" reactiontime="+66" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202663" lastname="COOPER" firstname="Isaac Alan" gender="M" birthdate="2004-01-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.43" eventid="3" heat="3" lane="2">
                  <MEETINFO date="2021-07-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.31" eventid="19" heat="6" lane="2">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="3" lane="1" heat="1" heatid="10103" swimtime="00:00:49.52" reactiontime="+59" points="929">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:23.78" />
                    <SPLIT distance="75" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:00:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="6" lane="2" heat="3" heatid="30003" swimtime="00:00:50.16" reactiontime="+57" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                    <SPLIT distance="75" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:00:50.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="7" lane="3" heat="1" heatid="10203" swimtime="00:00:50.01" reactiontime="+57" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:23.95" />
                    <SPLIT distance="75" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="2" lane="4" heat="1" heatid="10119" swimtime="00:00:22.73" reactiontime="+53" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.06" />
                    <SPLIT distance="50" swimtime="00:00:22.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="2" lane="2" heat="6" heatid="60019" swimtime="00:00:22.79" reactiontime="+59" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.18" />
                    <SPLIT distance="50" swimtime="00:00:22.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="1" lane="4" heat="1" heatid="10219" swimtime="00:00:22.52" reactiontime="+56" points="960">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.01" />
                    <SPLIT distance="50" swimtime="00:00:22.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163641" lastname="YONG" firstname="Joshua" gender="M" birthdate="2001-07-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.63" eventid="16" heat="7" lane="8">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="14" lane="8" heat="7" heatid="70016" swimtime="00:00:57.77" reactiontime="+74" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.44" />
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                    <SPLIT distance="75" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:00:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="10" lane="1" heat="1" heatid="10216" swimtime="00:00:57.34" reactiontime="+69" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="75" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:00:57.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191499" lastname="WILLIAMSON" firstname="Sam" gender="M" birthdate="1997-12-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.01" eventid="16" heat="8" lane="6">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.27" eventid="41" heat="8" lane="2">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="23" lane="6" heat="8" heatid="80016" swimtime="00:00:58.13" reactiontime="+65" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:42.49" />
                    <SPLIT distance="100" swimtime="00:00:58.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="13" lane="2" heat="8" heatid="80041" swimtime="00:00:26.42" reactiontime="+64" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="11" lane="1" heat="2" heatid="20241" swimtime="00:00:26.25" reactiontime="+64" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156743" lastname="TEMPLE" firstname="Matthew" gender="M" birthdate="1999-06-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.68" eventid="39" heat="7" lane="3">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.78" eventid="14" heat="10" lane="2">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.70" eventid="5" heat="10" lane="1">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="7" lane="1" heat="1" heatid="10139" swimtime="00:00:49.67" reactiontime="+62" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.94" />
                    <SPLIT distance="75" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:00:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="5" lane="3" heat="7" heatid="70039" swimtime="00:00:49.85" reactiontime="+65" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.70" />
                    <SPLIT distance="50" swimtime="00:00:23.22" />
                    <SPLIT distance="75" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:00:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="7" lane="3" heat="2" heatid="20239" swimtime="00:00:49.73" reactiontime="+65" points="886">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.36" />
                    <SPLIT distance="75" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:00:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="15" lane="2" heat="10" heatid="100014" swimtime="00:00:46.98" reactiontime="+63" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.71" />
                    <SPLIT distance="75" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:00:46.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="13" lane="8" heat="2" heatid="20214" swimtime="00:00:46.63" reactiontime="+62" points="889">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.64" />
                    <SPLIT distance="50" swimtime="00:00:22.50" />
                    <SPLIT distance="75" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:00:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="6" lane="1" heat="10" heatid="100005" swimtime="00:00:22.30" reactiontime="+62" points="927">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.26" />
                    <SPLIT distance="50" swimtime="00:00:22.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="12" lane="3" heat="1" heatid="10205" swimtime="00:00:22.37" reactiontime="+60" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.34" />
                    <SPLIT distance="50" swimtime="00:00:22.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202666" lastname="CHAMPION" firstname="Shaun" gender="M" birthdate="2000-03-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.31" eventid="39" heat="8" lane="1">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="13" lane="1" heat="8" heatid="80039" swimtime="00:00:50.54" reactiontime="+61" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.64" />
                    <SPLIT distance="50" swimtime="00:00:23.39" />
                    <SPLIT distance="75" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:00:50.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="13" lane="1" heat="2" heatid="20239" swimtime="00:00:50.56" reactiontime="+62" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.72" />
                    <SPLIT distance="50" swimtime="00:00:23.62" />
                    <SPLIT distance="75" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120880" lastname="CHALMERS" firstname="Kyle" gender="M" birthdate="1998-06-25">
              <ENTRIES>
                <ENTRY entrytime="00:00:44.84" eventid="14" heat="11" lane="4">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:40.82" eventid="44" heat="5" lane="4">
                  <MEETINFO date="2021-10-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:20.68" eventid="31" heat="10" lane="4">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="1" lane="3" heat="1" heatid="10114" swimtime="00:00:45.16" reactiontime="+67" points="978">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.63" />
                    <SPLIT distance="75" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:00:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="3" lane="4" heat="11" heatid="110014" swimtime="00:00:45.84" reactiontime="+70" points="935">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.41" />
                    <SPLIT distance="50" swimtime="00:00:22.04" />
                    <SPLIT distance="75" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:00:45.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="3" lane="5" heat="2" heatid="20214" swimtime="00:00:45.66" reactiontime="+67" points="947">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.29" />
                    <SPLIT distance="50" swimtime="00:00:21.93" />
                    <SPLIT distance="75" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="-1" lane="4" heat="5" heatid="50044" swimtime="NT" status="DNS" />
                <RESULT eventid="131" place="7" lane="6" heat="1" heatid="10131" swimtime="00:00:20.92" reactiontime="+68" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.18" />
                    <SPLIT distance="50" swimtime="00:00:20.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="9" lane="4" heat="10" heatid="100031" swimtime="00:00:21.09" reactiontime="+68" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.22" />
                    <SPLIT distance="50" swimtime="00:00:21.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="4" lane="6" heat="1" heatid="10231" swimtime="00:00:20.91" reactiontime="+67" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.12" />
                    <SPLIT distance="50" swimtime="00:00:20.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150388" lastname="SWINBURN" firstname="Stuart" gender="M" birthdate="2001-06-23">
              <ENTRIES>
                <ENTRY entrytime="00:14:47.96" eventid="10" heat="2" lane="2">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="10" lane="2" heat="2" heatid="20010" swimtime="00:14:51.00" reactiontime="+72" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                    <SPLIT distance="75" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:00:54.86" />
                    <SPLIT distance="125" swimtime="00:01:09.61" />
                    <SPLIT distance="150" swimtime="00:01:24.32" />
                    <SPLIT distance="175" swimtime="00:01:39.16" />
                    <SPLIT distance="200" swimtime="00:01:54.09" />
                    <SPLIT distance="225" swimtime="00:02:08.89" />
                    <SPLIT distance="250" swimtime="00:02:23.77" />
                    <SPLIT distance="275" swimtime="00:02:38.70" />
                    <SPLIT distance="300" swimtime="00:02:53.56" />
                    <SPLIT distance="325" swimtime="00:03:08.42" />
                    <SPLIT distance="350" swimtime="00:03:23.35" />
                    <SPLIT distance="375" swimtime="00:03:38.25" />
                    <SPLIT distance="400" swimtime="00:03:53.26" />
                    <SPLIT distance="425" swimtime="00:04:08.09" />
                    <SPLIT distance="450" swimtime="00:04:22.99" />
                    <SPLIT distance="475" swimtime="00:04:37.87" />
                    <SPLIT distance="500" swimtime="00:04:52.77" />
                    <SPLIT distance="525" swimtime="00:05:07.72" />
                    <SPLIT distance="550" swimtime="00:05:22.63" />
                    <SPLIT distance="575" swimtime="00:05:37.47" />
                    <SPLIT distance="600" swimtime="00:05:52.30" />
                    <SPLIT distance="625" swimtime="00:06:07.13" />
                    <SPLIT distance="650" swimtime="00:06:22.08" />
                    <SPLIT distance="675" swimtime="00:06:36.94" />
                    <SPLIT distance="700" swimtime="00:06:52.00" />
                    <SPLIT distance="725" swimtime="00:07:07.16" />
                    <SPLIT distance="750" swimtime="00:07:22.28" />
                    <SPLIT distance="775" swimtime="00:07:37.38" />
                    <SPLIT distance="800" swimtime="00:07:52.35" />
                    <SPLIT distance="825" swimtime="00:08:07.40" />
                    <SPLIT distance="850" swimtime="00:08:22.38" />
                    <SPLIT distance="875" swimtime="00:08:37.34" />
                    <SPLIT distance="900" swimtime="00:08:52.35" />
                    <SPLIT distance="925" swimtime="00:09:07.42" />
                    <SPLIT distance="950" swimtime="00:09:22.32" />
                    <SPLIT distance="975" swimtime="00:09:37.19" />
                    <SPLIT distance="1000" swimtime="00:09:52.25" />
                    <SPLIT distance="1025" swimtime="00:10:07.24" />
                    <SPLIT distance="1050" swimtime="00:10:22.36" />
                    <SPLIT distance="1075" swimtime="00:10:37.30" />
                    <SPLIT distance="1100" swimtime="00:10:52.34" />
                    <SPLIT distance="1125" swimtime="00:11:07.32" />
                    <SPLIT distance="1150" swimtime="00:11:22.35" />
                    <SPLIT distance="1175" swimtime="00:11:37.55" />
                    <SPLIT distance="1200" swimtime="00:11:52.55" />
                    <SPLIT distance="1225" swimtime="00:12:07.64" />
                    <SPLIT distance="1250" swimtime="00:12:22.68" />
                    <SPLIT distance="1275" swimtime="00:12:37.92" />
                    <SPLIT distance="1300" swimtime="00:12:52.97" />
                    <SPLIT distance="1325" swimtime="00:13:08.00" />
                    <SPLIT distance="1350" swimtime="00:13:23.01" />
                    <SPLIT distance="1375" swimtime="00:13:38.00" />
                    <SPLIT distance="1400" swimtime="00:13:53.11" />
                    <SPLIT distance="1425" swimtime="00:14:08.19" />
                    <SPLIT distance="1450" swimtime="00:14:23.07" />
                    <SPLIT distance="1475" swimtime="00:14:37.51" />
                    <SPLIT distance="1500" swimtime="00:14:51.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163630" lastname="HARTWELL" firstname="Ty" gender="M" birthdate="2001-01-10">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.28" eventid="46" heat="3" lane="2">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="11" lane="2" heat="3" heatid="30046" swimtime="00:01:51.95" reactiontime="+56" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:26.46" />
                    <SPLIT distance="75" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:00:55.14" />
                    <SPLIT distance="125" swimtime="00:01:09.17" />
                    <SPLIT distance="150" swimtime="00:01:23.41" />
                    <SPLIT distance="175" swimtime="00:01:37.97" />
                    <SPLIT distance="200" swimtime="00:01:51.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150360" lastname="SCHLICHT" firstname="David" gender="M" birthdate="1999-09-03">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.79" eventid="29" heat="5" lane="8">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="00:04:01.44" eventid="37" heat="3" lane="3">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="29" place="16" lane="8" heat="5" heatid="50029" swimtime="00:02:06.72" reactiontime="+66" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="75" swimtime="00:00:44.57" />
                    <SPLIT distance="100" swimtime="00:01:00.67" />
                    <SPLIT distance="125" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:33.37" />
                    <SPLIT distance="175" swimtime="00:01:50.06" />
                    <SPLIT distance="200" swimtime="00:02:06.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="7" lane="2" heat="1" heatid="10137" swimtime="00:04:04.33" reactiontime="+65" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                    <SPLIT distance="75" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:00:55.72" />
                    <SPLIT distance="125" swimtime="00:01:11.84" />
                    <SPLIT distance="150" swimtime="00:01:27.44" />
                    <SPLIT distance="175" swimtime="00:01:43.10" />
                    <SPLIT distance="200" swimtime="00:01:58.72" />
                    <SPLIT distance="225" swimtime="00:02:15.86" />
                    <SPLIT distance="250" swimtime="00:02:33.01" />
                    <SPLIT distance="275" swimtime="00:02:50.37" />
                    <SPLIT distance="300" swimtime="00:03:07.74" />
                    <SPLIT distance="325" swimtime="00:03:22.39" />
                    <SPLIT distance="350" swimtime="00:03:36.52" />
                    <SPLIT distance="375" swimtime="00:03:50.62" />
                    <SPLIT distance="400" swimtime="00:04:04.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="5" lane="3" heat="3" heatid="30037" swimtime="00:04:02.85" reactiontime="+63" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                    <SPLIT distance="75" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:00:55.58" />
                    <SPLIT distance="125" swimtime="00:01:11.38" />
                    <SPLIT distance="150" swimtime="00:01:26.71" />
                    <SPLIT distance="175" swimtime="00:01:42.18" />
                    <SPLIT distance="200" swimtime="00:01:57.45" />
                    <SPLIT distance="225" swimtime="00:02:14.22" />
                    <SPLIT distance="250" swimtime="00:02:31.11" />
                    <SPLIT distance="275" swimtime="00:02:48.32" />
                    <SPLIT distance="300" swimtime="00:03:05.71" />
                    <SPLIT distance="325" swimtime="00:03:20.45" />
                    <SPLIT distance="350" swimtime="00:03:34.77" />
                    <SPLIT distance="375" swimtime="00:03:49.05" />
                    <SPLIT distance="400" swimtime="00:04:02.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163637" lastname="NEILL" firstname="Thomas" gender="M" birthdate="2002-06-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.56" eventid="44" heat="4" lane="6">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:03:38.24" eventid="24" heat="4" lane="6">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="144" place="5" lane="1" heat="1" heatid="10144" swimtime="00:01:41.55" reactiontime="+65" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.25" />
                    <SPLIT distance="50" swimtime="00:00:23.77" />
                    <SPLIT distance="75" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:00:49.49" />
                    <SPLIT distance="125" swimtime="00:01:02.49" />
                    <SPLIT distance="150" swimtime="00:01:15.80" />
                    <SPLIT distance="175" swimtime="00:01:28.98" />
                    <SPLIT distance="200" swimtime="00:01:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="7" lane="6" heat="4" heatid="40044" swimtime="00:01:42.38" reactiontime="+66" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:24.09" />
                    <SPLIT distance="75" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:00:50.06" />
                    <SPLIT distance="125" swimtime="00:01:03.21" />
                    <SPLIT distance="150" swimtime="00:01:16.50" />
                    <SPLIT distance="175" swimtime="00:01:29.67" />
                    <SPLIT distance="200" swimtime="00:01:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="124" place="2" lane="2" heat="1" heatid="10124" swimtime="00:03:35.05" reactiontime="+67" points="961">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                    <SPLIT distance="75" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:00:51.65" />
                    <SPLIT distance="125" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:18.76" />
                    <SPLIT distance="175" swimtime="00:01:32.31" />
                    <SPLIT distance="200" swimtime="00:01:45.99" />
                    <SPLIT distance="225" swimtime="00:01:59.63" />
                    <SPLIT distance="250" swimtime="00:02:13.41" />
                    <SPLIT distance="275" swimtime="00:02:27.07" />
                    <SPLIT distance="300" swimtime="00:02:40.77" />
                    <SPLIT distance="325" swimtime="00:02:54.43" />
                    <SPLIT distance="350" swimtime="00:03:08.16" />
                    <SPLIT distance="375" swimtime="00:03:21.89" />
                    <SPLIT distance="400" swimtime="00:03:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="5" lane="6" heat="4" heatid="40024" swimtime="00:03:38.23" reactiontime="+66" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                    <SPLIT distance="50" swimtime="00:00:25.17" />
                    <SPLIT distance="75" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:00:52.79" />
                    <SPLIT distance="125" swimtime="00:01:06.49" />
                    <SPLIT distance="150" swimtime="00:01:20.49" />
                    <SPLIT distance="175" swimtime="00:01:34.59" />
                    <SPLIT distance="200" swimtime="00:01:48.59" />
                    <SPLIT distance="225" swimtime="00:02:02.57" />
                    <SPLIT distance="250" swimtime="00:02:16.63" />
                    <SPLIT distance="275" swimtime="00:02:30.35" />
                    <SPLIT distance="300" swimtime="00:02:44.11" />
                    <SPLIT distance="325" swimtime="00:02:57.85" />
                    <SPLIT distance="350" swimtime="00:03:11.58" />
                    <SPLIT distance="375" swimtime="00:03:25.15" />
                    <SPLIT distance="400" swimtime="00:03:38.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120888" lastname="LEWIS" firstname="Clyde" gender="M" birthdate="1997-09-25">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.01" eventid="7" heat="5" lane="6">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:52.57" eventid="23" heat="3" lane="2">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="107" place="7" lane="7" heat="1" heatid="10107" swimtime="00:01:53.19" reactiontime="+72" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.19" />
                    <SPLIT distance="50" swimtime="00:00:24.66" />
                    <SPLIT distance="75" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:00:52.64" />
                    <SPLIT distance="125" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:26.16" />
                    <SPLIT distance="175" swimtime="00:01:40.39" />
                    <SPLIT distance="200" swimtime="00:01:53.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="6" lane="6" heat="5" heatid="50007" swimtime="00:01:52.83" reactiontime="+68" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.07" />
                    <SPLIT distance="50" swimtime="00:00:24.50" />
                    <SPLIT distance="75" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:00:52.58" />
                    <SPLIT distance="125" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:25.63" />
                    <SPLIT distance="175" swimtime="00:01:39.83" />
                    <SPLIT distance="200" swimtime="00:01:52.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="19" lane="2" heat="3" heatid="30023" swimtime="00:00:52.82" reactiontime="+68" points="812">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.65" />
                    <SPLIT distance="50" swimtime="00:00:23.99" />
                    <SPLIT distance="75" swimtime="00:00:39.51" />
                    <SPLIT distance="100" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173960" lastname="LEE" firstname="Se-Bom" gender="M" birthdate="2001-06-12">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.83" eventid="7" heat="5" lane="2">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="12" lane="2" heat="5" heatid="50007" swimtime="00:01:53.71" reactiontime="+63" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:24.66" />
                    <SPLIT distance="75" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:00:52.60" />
                    <SPLIT distance="125" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:26.04" />
                    <SPLIT distance="175" swimtime="00:01:40.40" />
                    <SPLIT distance="200" swimtime="00:01:53.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110896" lastname="HORTON" firstname="Mack" gender="M" birthdate="1996-04-25">
              <ENTRIES>
                <ENTRY entrytime="00:03:37.94" eventid="24" heat="4" lane="3">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:07:39.71" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="124" place="6" lane="6" heat="1" heatid="10124" swimtime="00:03:37.94" reactiontime="+71" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                    <SPLIT distance="75" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:00:52.62" />
                    <SPLIT distance="125" swimtime="00:01:06.38" />
                    <SPLIT distance="150" swimtime="00:01:20.16" />
                    <SPLIT distance="175" swimtime="00:01:34.00" />
                    <SPLIT distance="200" swimtime="00:01:48.00" />
                    <SPLIT distance="225" swimtime="00:02:01.77" />
                    <SPLIT distance="250" swimtime="00:02:15.85" />
                    <SPLIT distance="275" swimtime="00:02:29.73" />
                    <SPLIT distance="300" swimtime="00:02:43.96" />
                    <SPLIT distance="325" swimtime="00:02:57.57" />
                    <SPLIT distance="350" swimtime="00:03:11.40" />
                    <SPLIT distance="375" swimtime="00:03:25.03" />
                    <SPLIT distance="400" swimtime="00:03:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="4" lane="3" heat="4" heatid="40024" swimtime="00:03:38.09" reactiontime="+72" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:25.39" />
                    <SPLIT distance="75" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:00:53.11" />
                    <SPLIT distance="125" swimtime="00:01:06.79" />
                    <SPLIT distance="150" swimtime="00:01:20.87" />
                    <SPLIT distance="175" swimtime="00:01:34.73" />
                    <SPLIT distance="200" swimtime="00:01:48.63" />
                    <SPLIT distance="225" swimtime="00:02:02.35" />
                    <SPLIT distance="250" swimtime="00:02:16.30" />
                    <SPLIT distance="275" swimtime="00:02:30.18" />
                    <SPLIT distance="300" swimtime="00:02:44.12" />
                    <SPLIT distance="325" swimtime="00:02:57.86" />
                    <SPLIT distance="350" swimtime="00:03:11.68" />
                    <SPLIT distance="375" swimtime="00:03:25.36" />
                    <SPLIT distance="400" swimtime="00:03:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="9" lane="7" heat="5" heatid="30142" swimtime="00:07:40.64" reactiontime="+75" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                    <SPLIT distance="75" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:00:55.17" />
                    <SPLIT distance="125" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:23.72" />
                    <SPLIT distance="175" swimtime="00:01:37.69" />
                    <SPLIT distance="200" swimtime="00:01:51.99" />
                    <SPLIT distance="225" swimtime="00:02:06.11" />
                    <SPLIT distance="250" swimtime="00:02:20.60" />
                    <SPLIT distance="275" swimtime="00:02:34.83" />
                    <SPLIT distance="300" swimtime="00:02:49.28" />
                    <SPLIT distance="325" swimtime="00:03:03.43" />
                    <SPLIT distance="350" swimtime="00:03:17.97" />
                    <SPLIT distance="375" swimtime="00:03:32.28" />
                    <SPLIT distance="400" swimtime="00:03:46.86" />
                    <SPLIT distance="425" swimtime="00:04:01.18" />
                    <SPLIT distance="450" swimtime="00:04:15.74" />
                    <SPLIT distance="475" swimtime="00:04:30.02" />
                    <SPLIT distance="500" swimtime="00:04:44.52" />
                    <SPLIT distance="525" swimtime="00:04:58.83" />
                    <SPLIT distance="550" swimtime="00:05:13.47" />
                    <SPLIT distance="575" swimtime="00:05:27.91" />
                    <SPLIT distance="600" swimtime="00:05:42.68" />
                    <SPLIT distance="625" swimtime="00:05:57.35" />
                    <SPLIT distance="650" swimtime="00:06:12.24" />
                    <SPLIT distance="675" swimtime="00:06:27.13" />
                    <SPLIT distance="700" swimtime="00:06:42.10" />
                    <SPLIT distance="725" swimtime="00:06:56.96" />
                    <SPLIT distance="750" swimtime="00:07:11.96" />
                    <SPLIT distance="775" swimtime="00:07:26.65" />
                    <SPLIT distance="800" swimtime="00:07:40.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202654" lastname="SMITH" firstname="Brendon Peter" gender="M" birthdate="2000-07-04">
              <ENTRIES>
                <ENTRY entrytime="00:03:59.33" eventid="37" heat="3" lane="5">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="37" place="-1" lane="5" heat="3" heatid="30037" swimtime="00:04:02.22" status="DSQ" reactiontime="+72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120878" lastname="BELL" firstname="Grayson" gender="M" birthdate="1997-03-21">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:26.45" eventid="41" heat="7" lane="7">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.36" eventid="31" heat="11" lane="1">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="11" lane="7" heat="7" heatid="70041" swimtime="00:00:26.37" reactiontime="+62" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:26.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="10" lane="7" heat="2" heatid="20241" swimtime="00:00:26.24" reactiontime="+62" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="25" lane="1" heat="11" heatid="110031" swimtime="00:00:21.42" reactiontime="+61" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:21.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130172" lastname="MCKEOWN" firstname="Kaylee" gender="F" birthdate="2001-07-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.81" eventid="2" heat="5" lane="5">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:01:59.48" eventid="45" heat="5" lane="4">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.63" eventid="6" heat="3" lane="5">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:26.32" eventid="18" heat="6" lane="6">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="1" lane="7" heat="1" heatid="10102" swimtime="00:00:55.49" reactiontime="+55" points="967">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.01" />
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                    <SPLIT distance="75" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:00:55.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="12" lane="5" heat="5" heatid="50002" swimtime="00:00:57.11" reactiontime="+55" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:42.66" />
                    <SPLIT distance="100" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="6" lane="7" heat="1" heatid="10202" swimtime="00:00:56.35" reactiontime="+54" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="1" lane="5" heat="1" heatid="10145" swimtime="00:01:59.26" reactiontime="+56" points="991">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:00:58.26" />
                    <SPLIT distance="125" swimtime="00:01:13.41" />
                    <SPLIT distance="150" swimtime="00:01:28.92" />
                    <SPLIT distance="175" swimtime="00:01:44.26" />
                    <SPLIT distance="200" swimtime="00:01:59.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="2" lane="4" heat="5" heatid="50045" swimtime="00:02:02.32" reactiontime="+58" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="75" swimtime="00:00:44.18" />
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="125" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:31.08" />
                    <SPLIT distance="175" swimtime="00:01:46.90" />
                    <SPLIT distance="200" swimtime="00:02:02.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106" place="3" lane="6" heat="1" heatid="10106" swimtime="00:02:03.57" reactiontime="+66" points="959">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                    <SPLIT distance="75" swimtime="00:00:42.86" />
                    <SPLIT distance="100" swimtime="00:00:57.66" />
                    <SPLIT distance="125" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:33.88" />
                    <SPLIT distance="175" swimtime="00:01:49.54" />
                    <SPLIT distance="200" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="4" lane="5" heat="3" heatid="30006" swimtime="00:02:06.07" reactiontime="+68" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="75" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:00:58.90" />
                    <SPLIT distance="125" swimtime="00:01:16.92" />
                    <SPLIT distance="150" swimtime="00:01:35.54" />
                    <SPLIT distance="175" swimtime="00:01:51.41" />
                    <SPLIT distance="200" swimtime="00:02:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="10" lane="6" heat="6" heatid="60018" swimtime="00:00:26.24" reactiontime="+56" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="9" lane="2" heat="1" heatid="10218" swimtime="00:00:26.09" reactiontime="+55" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.85" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163620" lastname="O'CALLAGHAN" firstname="Mollie" gender="F" birthdate="2004-04-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.02" eventid="2" heat="6" lane="3">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:26.52" eventid="18" heat="7" lane="7">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="2" lane="4" heat="1" heatid="10102" swimtime="00:00:55.62" reactiontime="+55" points="961">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                    <SPLIT distance="75" swimtime="00:00:41.12" />
                    <SPLIT distance="100" swimtime="00:00:55.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="3" lane="3" heat="6" heatid="60002" swimtime="00:00:56.35" reactiontime="+55" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                    <SPLIT distance="75" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="1" lane="5" heat="2" heatid="20202" swimtime="00:00:55.80" reactiontime="+53" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="75" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:00:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="3" lane="3" heat="1" heatid="10118" swimtime="00:00:25.61" reactiontime="+57" points="960">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="3" lane="7" heat="7" heatid="70018" swimtime="00:00:25.99" reactiontime="+56" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="3" lane="5" heat="2" heatid="20218" swimtime="00:00:25.69" reactiontime="+55" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129244" lastname="STRAUCH" firstname="Jenna" gender="F" birthdate="1997-03-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.20" eventid="15" heat="6" lane="7">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.94" eventid="28" heat="4" lane="3">
                  <MEETINFO date="2021-09-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:30.19" eventid="40" heat="5" lane="7">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="17" lane="7" heat="6" heatid="60015" swimtime="00:01:05.30" reactiontime="+71" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="75" swimtime="00:00:47.55" />
                    <SPLIT distance="100" swimtime="00:01:05.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="128" place="4" lane="7" heat="1" heatid="10128" swimtime="00:02:18.87" reactiontime="+71" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.50" />
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="75" swimtime="00:00:49.22" />
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                    <SPLIT distance="125" swimtime="00:01:24.74" />
                    <SPLIT distance="150" swimtime="00:01:42.62" />
                    <SPLIT distance="175" swimtime="00:02:00.55" />
                    <SPLIT distance="200" swimtime="00:02:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="6" lane="3" heat="4" heatid="40028" swimtime="00:02:19.75" reactiontime="+69" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="75" swimtime="00:00:49.20" />
                    <SPLIT distance="100" swimtime="00:01:06.74" />
                    <SPLIT distance="125" swimtime="00:01:24.32" />
                    <SPLIT distance="150" swimtime="00:01:42.27" />
                    <SPLIT distance="175" swimtime="00:02:00.77" />
                    <SPLIT distance="200" swimtime="00:02:19.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="-1" lane="7" heat="5" heatid="50040" swimtime="00:00:30.26" status="DSQ" reactiontime="+70" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150358" lastname="HODGES" firstname="Chelsea" gender="F" birthdate="2001-06-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.78" eventid="15" heat="7" lane="6">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:29.91" eventid="40" heat="7" lane="2">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="26" lane="6" heat="7" heatid="70015" swimtime="00:01:06.29" reactiontime="+71" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.09" />
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="75" swimtime="00:00:48.22" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="11" lane="2" heat="7" heatid="70040" swimtime="00:00:29.84" reactiontime="+65" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="9" lane="7" heat="2" heatid="20240" swimtime="00:00:29.85" reactiontime="+68" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172303" lastname="CASTELLUZZO" firstname="Brittany" gender="F" birthdate="2000-11-26">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.18" eventid="38" heat="2" lane="2">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="16" lane="2" heat="2" heatid="20038" swimtime="00:00:57.85" reactiontime="+60" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:00:57.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="338" place="17" lane="4" heat="1" heatid="10338" swimtime="00:00:57.76" reactiontime="+61" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                    <SPLIT distance="75" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:00:57.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202753" lastname="PERKINS" firstname="Alexandria" gender="F" birthdate="2000-07-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.89" eventid="38" heat="3" lane="6">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.52" eventid="4" heat="4" lane="2">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="138" place="6" lane="2" heat="1" heatid="10138" swimtime="00:00:56.34" reactiontime="+70" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.03" />
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                    <SPLIT distance="75" swimtime="00:00:41.00" />
                    <SPLIT distance="100" swimtime="00:00:56.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="3" lane="6" heat="3" heatid="30038" swimtime="00:00:56.46" reactiontime="+69" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                    <SPLIT distance="75" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:00:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="6" lane="5" heat="2" heatid="20238" swimtime="00:00:56.39" reactiontime="+68" points="907">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:26.37" />
                    <SPLIT distance="75" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:00:56.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="16" lane="2" heat="4" heatid="40004" swimtime="00:00:25.65" reactiontime="+74" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:25.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="15" lane="8" heat="1" heatid="10204" swimtime="00:00:25.60" reactiontime="+72" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100650" lastname="MCKEON" firstname="Emma" gender="F" birthdate="1994-05-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:50.58" eventid="13" heat="9" lane="4">
                  <MEETINFO date="2021-10-09" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:23.50" eventid="30" heat="7" lane="4">
                  <MEETINFO date="2021-10-07" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="1" lane="4" heat="1" heatid="10113" swimtime="00:00:50.77" reactiontime="+72" points="969">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:24.41" />
                    <SPLIT distance="75" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:00:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="2" lane="4" heat="9" heatid="90013" swimtime="00:00:52.23" reactiontime="+74" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:24.88" />
                    <SPLIT distance="75" swimtime="00:00:38.56" />
                    <SPLIT distance="100" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="1" lane="5" heat="2" heatid="20213" swimtime="00:00:51.28" reactiontime="+74" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:24.62" />
                    <SPLIT distance="75" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="1" lane="5" heat="1" heatid="10130" swimtime="00:00:23.04" reactiontime="+70" points="985">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:23.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="6" lane="4" heat="7" heatid="70030" swimtime="00:00:23.93" reactiontime="+75" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.64" />
                    <SPLIT distance="50" swimtime="00:00:23.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="2" lane="3" heat="1" heatid="10230" swimtime="00:00:23.51" reactiontime="+74" points="927">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:23.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105256" lastname="WILSON" firstname="Madison" gender="F" birthdate="1994-05-31">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:51.40" eventid="13" heat="7" lane="4">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.23" eventid="43" heat="3" lane="4">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="4" lane="3" heat="1" heatid="10113" swimtime="00:00:51.70" reactiontime="+69" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                    <SPLIT distance="75" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:00:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="5" lane="4" heat="7" heatid="70013" swimtime="00:00:52.43" reactiontime="+67" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:25.59" />
                    <SPLIT distance="75" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:00:52.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="3" lane="3" heat="2" heatid="20213" swimtime="00:00:51.82" reactiontime="+69" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:00:51.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="143" place="8" lane="8" heat="1" heatid="10143" swimtime="00:01:53.39" reactiontime="+69" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.48" />
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                    <SPLIT distance="75" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:00:55.17" />
                    <SPLIT distance="125" swimtime="00:01:09.80" />
                    <SPLIT distance="150" swimtime="00:01:24.46" />
                    <SPLIT distance="175" swimtime="00:01:39.07" />
                    <SPLIT distance="200" swimtime="00:01:53.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="8" lane="4" heat="3" heatid="30043" swimtime="00:01:54.18" reactiontime="+68" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="75" swimtime="00:00:41.02" />
                    <SPLIT distance="100" swimtime="00:00:55.46" />
                    <SPLIT distance="125" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:24.81" />
                    <SPLIT distance="175" swimtime="00:01:39.70" />
                    <SPLIT distance="200" swimtime="00:01:54.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120863" lastname="ATHERTON" firstname="Minna" gender="F" birthdate="2000-05-17">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.40" eventid="45" heat="3" lane="4">
                  <MEETINFO date="2021-09-11" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="12" lane="4" heat="3" heatid="30045" swimtime="00:02:05.05" reactiontime="+58" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="75" swimtime="00:00:44.43" />
                    <SPLIT distance="100" swimtime="00:01:00.34" />
                    <SPLIT distance="125" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:32.53" />
                    <SPLIT distance="175" swimtime="00:01:49.14" />
                    <SPLIT distance="200" swimtime="00:02:05.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202759" lastname="SMITH" firstname="Mikayla Maree" gender="F" birthdate="1998-10-06">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.97" eventid="28" heat="5" lane="1">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="11" lane="1" heat="5" heatid="50028" swimtime="00:02:20.67" reactiontime="+63" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="75" swimtime="00:00:49.07" />
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                    <SPLIT distance="125" swimtime="00:01:25.24" />
                    <SPLIT distance="150" swimtime="00:01:43.52" />
                    <SPLIT distance="175" swimtime="00:02:01.78" />
                    <SPLIT distance="200" swimtime="00:02:20.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161731" lastname="TAYLOR" firstname="Laura" gender="F" birthdate="1999-09-10">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.91" eventid="20" heat="2" lane="6">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="9" lane="6" heat="2" heatid="20020" swimtime="00:02:05.94" reactiontime="+71" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                    <SPLIT distance="75" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:00.81" />
                    <SPLIT distance="125" swimtime="00:01:17.14" />
                    <SPLIT distance="150" swimtime="00:01:33.35" />
                    <SPLIT distance="175" swimtime="00:01:49.67" />
                    <SPLIT distance="200" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163613" lastname="DEKKERS" firstname="Elizabeth" gender="F" birthdate="2004-05-06">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.65" eventid="20" heat="4" lane="6">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="120" place="3" lane="1" heat="1" heatid="10120" swimtime="00:02:03.94" reactiontime="+70" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="75" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:00:59.77" />
                    <SPLIT distance="125" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:31.48" />
                    <SPLIT distance="175" swimtime="00:01:47.61" />
                    <SPLIT distance="200" swimtime="00:02:03.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="7" lane="6" heat="4" heatid="40020" swimtime="00:02:05.41" reactiontime="+70" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="75" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="125" swimtime="00:01:16.66" />
                    <SPLIT distance="150" swimtime="00:01:32.55" />
                    <SPLIT distance="175" swimtime="00:01:48.84" />
                    <SPLIT distance="200" swimtime="00:02:05.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="111247" lastname="NEALE" firstname="Leah" gender="F" birthdate="1995-08-01">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.22" eventid="43" heat="3" lane="5">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:04:01.28" eventid="1" heat="3" lane="3">
                  <MEETINFO date="2021-09-09" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="143" place="6" lane="7" heat="1" heatid="10143" swimtime="00:01:52.84" reactiontime="+68" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                    <SPLIT distance="75" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:00:55.07" />
                    <SPLIT distance="125" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:24.06" />
                    <SPLIT distance="175" swimtime="00:01:38.63" />
                    <SPLIT distance="200" swimtime="00:01:52.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="6" lane="5" heat="3" heatid="30043" swimtime="00:01:54.05" reactiontime="+68" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                    <SPLIT distance="75" swimtime="00:00:41.27" />
                    <SPLIT distance="100" swimtime="00:00:55.78" />
                    <SPLIT distance="125" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:24.94" />
                    <SPLIT distance="175" swimtime="00:01:39.77" />
                    <SPLIT distance="200" swimtime="00:01:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="101" place="8" lane="8" heat="1" heatid="10101" swimtime="00:04:03.45" reactiontime="+70" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="75" swimtime="00:00:42.51" />
                    <SPLIT distance="100" swimtime="00:00:57.85" />
                    <SPLIT distance="125" swimtime="00:01:12.97" />
                    <SPLIT distance="150" swimtime="00:01:28.68" />
                    <SPLIT distance="175" swimtime="00:01:44.31" />
                    <SPLIT distance="200" swimtime="00:01:59.94" />
                    <SPLIT distance="225" swimtime="00:02:15.48" />
                    <SPLIT distance="250" swimtime="00:02:31.13" />
                    <SPLIT distance="275" swimtime="00:02:46.75" />
                    <SPLIT distance="300" swimtime="00:03:02.37" />
                    <SPLIT distance="325" swimtime="00:03:17.92" />
                    <SPLIT distance="350" swimtime="00:03:33.26" />
                    <SPLIT distance="375" swimtime="00:03:48.77" />
                    <SPLIT distance="400" swimtime="00:04:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="8" lane="3" heat="3" heatid="30001" swimtime="00:04:02.30" reactiontime="+70" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="75" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:00:58.73" />
                    <SPLIT distance="125" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:29.53" />
                    <SPLIT distance="175" swimtime="00:01:44.78" />
                    <SPLIT distance="200" swimtime="00:02:00.15" />
                    <SPLIT distance="225" swimtime="00:02:15.55" />
                    <SPLIT distance="250" swimtime="00:02:30.87" />
                    <SPLIT distance="275" swimtime="00:02:46.16" />
                    <SPLIT distance="300" swimtime="00:03:01.49" />
                    <SPLIT distance="325" swimtime="00:03:16.82" />
                    <SPLIT distance="350" swimtime="00:03:32.37" />
                    <SPLIT distance="375" swimtime="00:03:47.83" />
                    <SPLIT distance="400" swimtime="00:04:02.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213818" lastname="HARDY" firstname="Kayla" gender="F" birthdate="2003-04-09">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.69" eventid="6" heat="5" lane="7">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="00:04:32.84" eventid="36" heat="3" lane="2">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.67" eventid="22" heat="2" lane="7">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="12" lane="7" heat="5" heatid="50006" swimtime="00:02:08.11" reactiontime="+68" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:43.82" />
                    <SPLIT distance="100" swimtime="00:00:59.69" />
                    <SPLIT distance="125" swimtime="00:01:18.20" />
                    <SPLIT distance="150" swimtime="00:01:37.04" />
                    <SPLIT distance="175" swimtime="00:01:53.16" />
                    <SPLIT distance="200" swimtime="00:02:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="10" lane="2" heat="3" heatid="30036" swimtime="00:04:34.77" reactiontime="+68" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.57" />
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="75" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:00.91" />
                    <SPLIT distance="125" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:01:35.13" />
                    <SPLIT distance="175" swimtime="00:01:52.32" />
                    <SPLIT distance="200" swimtime="00:02:09.43" />
                    <SPLIT distance="225" swimtime="00:02:28.50" />
                    <SPLIT distance="250" swimtime="00:02:48.11" />
                    <SPLIT distance="275" swimtime="00:03:07.98" />
                    <SPLIT distance="300" swimtime="00:03:28.20" />
                    <SPLIT distance="325" swimtime="00:03:45.29" />
                    <SPLIT distance="350" swimtime="00:04:01.58" />
                    <SPLIT distance="375" swimtime="00:04:18.27" />
                    <SPLIT distance="400" swimtime="00:04:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="16" lane="7" heat="2" heatid="20022" swimtime="00:01:00.16" reactiontime="+67" points="828">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                    <SPLIT distance="75" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="15" lane="8" heat="1" heatid="10222" swimtime="00:00:59.75" reactiontime="+69" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                    <SPLIT distance="75" swimtime="00:00:44.90" />
                    <SPLIT distance="100" swimtime="00:00:59.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150371" lastname="PALLISTER" firstname="Lani" gender="F" birthdate="2002-06-06">
              <ENTRIES>
                <ENTRY entrytime="00:03:56.74" eventid="1" heat="3" lane="4">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:08:07.37" eventid="12" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="00:15:24.63" eventid="33" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="101" place="1" lane="5" heat="1" heatid="10101" swimtime="00:03:55.04" reactiontime="+67" points="985">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.69" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:00:56.81" />
                    <SPLIT distance="125" swimtime="00:01:11.68" />
                    <SPLIT distance="150" swimtime="00:01:26.74" />
                    <SPLIT distance="175" swimtime="00:01:41.79" />
                    <SPLIT distance="200" swimtime="00:01:56.81" />
                    <SPLIT distance="225" swimtime="00:02:11.63" />
                    <SPLIT distance="250" swimtime="00:02:26.76" />
                    <SPLIT distance="275" swimtime="00:02:41.63" />
                    <SPLIT distance="300" swimtime="00:02:56.47" />
                    <SPLIT distance="325" swimtime="00:03:11.13" />
                    <SPLIT distance="350" swimtime="00:03:25.94" />
                    <SPLIT distance="375" swimtime="00:03:40.68" />
                    <SPLIT distance="400" swimtime="00:03:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="2" lane="4" heat="3" heatid="30001" swimtime="00:03:59.50" reactiontime="+69" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="75" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:00:56.59" />
                    <SPLIT distance="125" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:26.56" />
                    <SPLIT distance="175" swimtime="00:01:41.84" />
                    <SPLIT distance="200" swimtime="00:01:56.88" />
                    <SPLIT distance="225" swimtime="00:02:12.21" />
                    <SPLIT distance="250" swimtime="00:02:27.41" />
                    <SPLIT distance="275" swimtime="00:02:42.79" />
                    <SPLIT distance="300" swimtime="00:02:58.24" />
                    <SPLIT distance="325" swimtime="00:03:13.69" />
                    <SPLIT distance="350" swimtime="00:03:29.33" />
                    <SPLIT distance="375" swimtime="00:03:44.82" />
                    <SPLIT distance="400" swimtime="00:03:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="1" lane="4" heat="5" heatid="30112" swimtime="00:08:04.07" reactiontime="+69" points="970">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="75" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:00:57.72" />
                    <SPLIT distance="125" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:27.76" />
                    <SPLIT distance="175" swimtime="00:01:42.96" />
                    <SPLIT distance="200" swimtime="00:01:57.96" />
                    <SPLIT distance="225" swimtime="00:02:13.40" />
                    <SPLIT distance="250" swimtime="00:02:28.48" />
                    <SPLIT distance="275" swimtime="00:02:43.70" />
                    <SPLIT distance="300" swimtime="00:02:59.04" />
                    <SPLIT distance="325" swimtime="00:03:14.37" />
                    <SPLIT distance="350" swimtime="00:03:29.76" />
                    <SPLIT distance="375" swimtime="00:03:44.94" />
                    <SPLIT distance="400" swimtime="00:04:00.23" />
                    <SPLIT distance="425" swimtime="00:04:15.52" />
                    <SPLIT distance="450" swimtime="00:04:30.65" />
                    <SPLIT distance="475" swimtime="00:04:45.82" />
                    <SPLIT distance="500" swimtime="00:05:01.16" />
                    <SPLIT distance="525" swimtime="00:05:16.43" />
                    <SPLIT distance="550" swimtime="00:05:31.74" />
                    <SPLIT distance="575" swimtime="00:05:47.19" />
                    <SPLIT distance="600" swimtime="00:06:02.57" />
                    <SPLIT distance="625" swimtime="00:06:17.79" />
                    <SPLIT distance="650" swimtime="00:06:33.00" />
                    <SPLIT distance="675" swimtime="00:06:48.35" />
                    <SPLIT distance="700" swimtime="00:07:03.67" />
                    <SPLIT distance="725" swimtime="00:07:19.09" />
                    <SPLIT distance="750" swimtime="00:07:34.52" />
                    <SPLIT distance="775" swimtime="00:07:49.71" />
                    <SPLIT distance="800" swimtime="00:08:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="1" lane="4" heat="5" heatid="30133" swimtime="00:15:21.43" reactiontime="+63" points="988">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.83" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:42.57" />
                    <SPLIT distance="100" swimtime="00:00:57.65" />
                    <SPLIT distance="125" swimtime="00:01:12.94" />
                    <SPLIT distance="150" swimtime="00:01:28.25" />
                    <SPLIT distance="175" swimtime="00:01:43.79" />
                    <SPLIT distance="200" swimtime="00:01:59.11" />
                    <SPLIT distance="225" swimtime="00:02:14.50" />
                    <SPLIT distance="250" swimtime="00:02:29.83" />
                    <SPLIT distance="275" swimtime="00:02:45.25" />
                    <SPLIT distance="300" swimtime="00:03:00.44" />
                    <SPLIT distance="325" swimtime="00:03:15.72" />
                    <SPLIT distance="350" swimtime="00:03:30.96" />
                    <SPLIT distance="375" swimtime="00:03:46.17" />
                    <SPLIT distance="400" swimtime="00:04:01.43" />
                    <SPLIT distance="425" swimtime="00:04:16.67" />
                    <SPLIT distance="450" swimtime="00:04:31.90" />
                    <SPLIT distance="475" swimtime="00:04:47.35" />
                    <SPLIT distance="500" swimtime="00:05:02.79" />
                    <SPLIT distance="525" swimtime="00:05:18.39" />
                    <SPLIT distance="550" swimtime="00:05:33.73" />
                    <SPLIT distance="575" swimtime="00:05:49.20" />
                    <SPLIT distance="600" swimtime="00:06:04.55" />
                    <SPLIT distance="625" swimtime="00:06:20.16" />
                    <SPLIT distance="650" swimtime="00:06:35.53" />
                    <SPLIT distance="675" swimtime="00:06:51.17" />
                    <SPLIT distance="700" swimtime="00:07:06.72" />
                    <SPLIT distance="725" swimtime="00:07:22.24" />
                    <SPLIT distance="750" swimtime="00:07:37.76" />
                    <SPLIT distance="775" swimtime="00:07:53.20" />
                    <SPLIT distance="800" swimtime="00:08:08.66" />
                    <SPLIT distance="825" swimtime="00:08:23.98" />
                    <SPLIT distance="850" swimtime="00:08:39.38" />
                    <SPLIT distance="875" swimtime="00:08:54.81" />
                    <SPLIT distance="900" swimtime="00:09:10.40" />
                    <SPLIT distance="925" swimtime="00:09:25.88" />
                    <SPLIT distance="950" swimtime="00:09:41.45" />
                    <SPLIT distance="975" swimtime="00:09:56.88" />
                    <SPLIT distance="1000" swimtime="00:10:12.35" />
                    <SPLIT distance="1025" swimtime="00:10:27.66" />
                    <SPLIT distance="1050" swimtime="00:10:43.13" />
                    <SPLIT distance="1075" swimtime="00:10:58.53" />
                    <SPLIT distance="1100" swimtime="00:11:14.06" />
                    <SPLIT distance="1125" swimtime="00:11:29.47" />
                    <SPLIT distance="1150" swimtime="00:11:45.07" />
                    <SPLIT distance="1175" swimtime="00:12:00.53" />
                    <SPLIT distance="1200" swimtime="00:12:16.10" />
                    <SPLIT distance="1225" swimtime="00:12:31.70" />
                    <SPLIT distance="1250" swimtime="00:12:47.26" />
                    <SPLIT distance="1275" swimtime="00:13:02.73" />
                    <SPLIT distance="1300" swimtime="00:13:18.34" />
                    <SPLIT distance="1325" swimtime="00:13:33.98" />
                    <SPLIT distance="1350" swimtime="00:13:49.54" />
                    <SPLIT distance="1375" swimtime="00:14:05.06" />
                    <SPLIT distance="1400" swimtime="00:14:20.53" />
                    <SPLIT distance="1425" swimtime="00:14:36.14" />
                    <SPLIT distance="1450" swimtime="00:14:51.60" />
                    <SPLIT distance="1475" swimtime="00:15:06.89" />
                    <SPLIT distance="1500" swimtime="00:15:21.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202661" lastname="MUIR" firstname="Emilie" gender="F" birthdate="2003-04-10">
              <ENTRIES>
                <ENTRY entrytime="00:04:33.84" eventid="36" heat="3" lane="1">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="36" place="11" lane="1" heat="3" heatid="30036" swimtime="00:04:35.52" reactiontime="+81" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:29.33" />
                    <SPLIT distance="75" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:02.47" />
                    <SPLIT distance="125" swimtime="00:01:20.61" />
                    <SPLIT distance="150" swimtime="00:01:37.99" />
                    <SPLIT distance="175" swimtime="00:01:55.20" />
                    <SPLIT distance="200" swimtime="00:02:12.18" />
                    <SPLIT distance="225" swimtime="00:02:32.01" />
                    <SPLIT distance="250" swimtime="00:02:52.00" />
                    <SPLIT distance="275" swimtime="00:03:11.82" />
                    <SPLIT distance="300" swimtime="00:03:31.97" />
                    <SPLIT distance="325" swimtime="00:03:48.37" />
                    <SPLIT distance="350" swimtime="00:04:04.42" />
                    <SPLIT distance="375" swimtime="00:04:20.39" />
                    <SPLIT distance="400" swimtime="00:04:35.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="173958" lastname="HARRIS" firstname="Meg" gender="F" birthdate="2002-03-07">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:23.84" eventid="30" heat="6" lane="5">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="130" place="6" lane="7" heat="1" heatid="10130" swimtime="00:00:23.73" reactiontime="+69" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="2" lane="5" heat="6" heatid="60030" swimtime="00:00:23.77" reactiontime="+70" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.57" />
                    <SPLIT distance="50" swimtime="00:00:23.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="6" lane="4" heat="1" heatid="10230" swimtime="00:00:23.97" reactiontime="+69" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:23.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202768" lastname="PERKINS" firstname="Jamie Ann" gender="F" birthdate="2005-01-19">
              <ENTRIES>
                <ENTRY entrytime="00:08:30.03" eventid="12" heat="2" lane="7">
                  <MEETINFO date="2022-05-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="13" lane="7" heat="2" heatid="20012" swimtime="00:08:36.26" reactiontime="+78" points="800">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.78" />
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="75" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:00:59.94" />
                    <SPLIT distance="125" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:31.58" />
                    <SPLIT distance="175" swimtime="00:01:47.61" />
                    <SPLIT distance="200" swimtime="00:02:03.69" />
                    <SPLIT distance="225" swimtime="00:02:19.82" />
                    <SPLIT distance="250" swimtime="00:02:35.83" />
                    <SPLIT distance="275" swimtime="00:02:51.95" />
                    <SPLIT distance="300" swimtime="00:03:08.07" />
                    <SPLIT distance="325" swimtime="00:03:24.47" />
                    <SPLIT distance="350" swimtime="00:03:40.63" />
                    <SPLIT distance="375" swimtime="00:03:56.87" />
                    <SPLIT distance="400" swimtime="00:04:13.06" />
                    <SPLIT distance="425" swimtime="00:04:29.47" />
                    <SPLIT distance="450" swimtime="00:04:45.86" />
                    <SPLIT distance="475" swimtime="00:05:02.43" />
                    <SPLIT distance="500" swimtime="00:05:18.78" />
                    <SPLIT distance="525" swimtime="00:05:35.28" />
                    <SPLIT distance="550" swimtime="00:05:51.82" />
                    <SPLIT distance="575" swimtime="00:06:08.35" />
                    <SPLIT distance="600" swimtime="00:06:24.85" />
                    <SPLIT distance="625" swimtime="00:06:41.33" />
                    <SPLIT distance="650" swimtime="00:06:57.88" />
                    <SPLIT distance="675" swimtime="00:07:14.49" />
                    <SPLIT distance="700" swimtime="00:07:31.14" />
                    <SPLIT distance="725" swimtime="00:07:47.71" />
                    <SPLIT distance="750" swimtime="00:08:04.19" />
                    <SPLIT distance="775" swimtime="00:08:20.53" />
                    <SPLIT distance="800" swimtime="00:08:36.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163629" lastname="GRANT" firstname="Alexander" gender="M" birthdate="2001-01-24">
              <ENTRIES>
                <ENTRY entrytime="00:07:40.18" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="142" place="14" lane="1" heat="5" heatid="30142" swimtime="00:07:48.25" reactiontime="+73" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="75" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:00:55.98" />
                    <SPLIT distance="125" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:25.30" />
                    <SPLIT distance="175" swimtime="00:01:39.91" />
                    <SPLIT distance="200" swimtime="00:01:54.79" />
                    <SPLIT distance="225" swimtime="00:02:09.46" />
                    <SPLIT distance="250" swimtime="00:02:24.21" />
                    <SPLIT distance="275" swimtime="00:02:38.85" />
                    <SPLIT distance="300" swimtime="00:02:53.72" />
                    <SPLIT distance="325" swimtime="00:03:08.32" />
                    <SPLIT distance="350" swimtime="00:03:23.03" />
                    <SPLIT distance="375" swimtime="00:03:37.64" />
                    <SPLIT distance="400" swimtime="00:03:52.39" />
                    <SPLIT distance="425" swimtime="00:04:06.88" />
                    <SPLIT distance="450" swimtime="00:04:21.59" />
                    <SPLIT distance="475" swimtime="00:04:36.17" />
                    <SPLIT distance="500" swimtime="00:04:50.78" />
                    <SPLIT distance="525" swimtime="00:05:05.29" />
                    <SPLIT distance="550" swimtime="00:05:20.04" />
                    <SPLIT distance="575" swimtime="00:05:34.80" />
                    <SPLIT distance="600" swimtime="00:05:49.76" />
                    <SPLIT distance="625" swimtime="00:06:04.43" />
                    <SPLIT distance="650" swimtime="00:06:19.37" />
                    <SPLIT distance="675" swimtime="00:06:34.39" />
                    <SPLIT distance="700" swimtime="00:06:49.66" />
                    <SPLIT distance="725" swimtime="00:07:04.80" />
                    <SPLIT distance="750" swimtime="00:07:19.57" />
                    <SPLIT distance="775" swimtime="00:07:34.10" />
                    <SPLIT distance="800" swimtime="00:07:48.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202662" lastname="SOUTHAM" firstname="Flynn Zareb" gender="M" birthdate="2005-06-05" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Australia">
              <RESULTS>
                <RESULT eventid="109" place="2" lane="6" heat="1" swimtime="00:03:04.63" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.01" />
                    <SPLIT distance="50" swimtime="00:00:23.01" />
                    <SPLIT distance="75" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:00:47.04" />
                    <SPLIT distance="125" swimtime="00:00:57.25" />
                    <SPLIT distance="150" swimtime="00:01:09.10" />
                    <SPLIT distance="175" swimtime="00:01:21.23" />
                    <SPLIT distance="200" swimtime="00:01:33.10" />
                    <SPLIT distance="225" swimtime="00:01:43.39" />
                    <SPLIT distance="250" swimtime="00:01:55.19" />
                    <SPLIT distance="275" swimtime="00:02:07.48" />
                    <SPLIT distance="300" swimtime="00:02:19.65" />
                    <SPLIT distance="325" swimtime="00:02:29.49" />
                    <SPLIT distance="350" swimtime="00:02:40.91" />
                    <SPLIT distance="375" swimtime="00:02:52.81" />
                    <SPLIT distance="400" swimtime="00:03:04.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202662" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="156743" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="163637" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="120880" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="4" lane="3" heat="1" swimtime="00:03:07.02" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.75" />
                    <SPLIT distance="50" swimtime="00:00:22.61" />
                    <SPLIT distance="75" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:00:47.00" />
                    <SPLIT distance="125" swimtime="00:00:57.63" />
                    <SPLIT distance="150" swimtime="00:01:09.67" />
                    <SPLIT distance="175" swimtime="00:01:21.68" />
                    <SPLIT distance="200" swimtime="00:01:33.55" />
                    <SPLIT distance="225" swimtime="00:01:44.02" />
                    <SPLIT distance="250" swimtime="00:01:56.17" />
                    <SPLIT distance="275" swimtime="00:02:08.66" />
                    <SPLIT distance="300" swimtime="00:02:21.04" />
                    <SPLIT distance="325" swimtime="00:02:31.30" />
                    <SPLIT distance="350" swimtime="00:02:43.11" />
                    <SPLIT distance="375" swimtime="00:02:55.25" />
                    <SPLIT distance="400" swimtime="00:03:07.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="163637" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="202662" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="202666" reactiontime="+36" />
                    <RELAYPOSITION number="4" athleteid="156743" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Australia">
              <RESULTS>
                <RESULT eventid="148" place="1" lane="2" heat="1" swimtime="00:03:18.98" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                    <SPLIT distance="50" swimtime="00:00:23.73" />
                    <SPLIT distance="75" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:00:49.46" />
                    <SPLIT distance="125" swimtime="00:01:01.34" />
                    <SPLIT distance="150" swimtime="00:01:15.77" />
                    <SPLIT distance="175" swimtime="00:01:30.50" />
                    <SPLIT distance="200" swimtime="00:01:46.01" />
                    <SPLIT distance="225" swimtime="00:01:55.96" />
                    <SPLIT distance="250" swimtime="00:02:08.30" />
                    <SPLIT distance="275" swimtime="00:02:21.01" />
                    <SPLIT distance="300" swimtime="00:02:34.35" />
                    <SPLIT distance="325" swimtime="00:02:44.21" />
                    <SPLIT distance="350" swimtime="00:02:55.57" />
                    <SPLIT distance="375" swimtime="00:03:07.22" />
                    <SPLIT distance="400" swimtime="00:03:18.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202663" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="163641" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="156743" reactiontime="+7" />
                    <RELAYPOSITION number="4" athleteid="120880" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="5" lane="6" heat="3" swimtime="00:03:25.02" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:24.26" />
                    <SPLIT distance="75" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:00:50.42" />
                    <SPLIT distance="125" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:17.19" />
                    <SPLIT distance="175" swimtime="00:01:32.32" />
                    <SPLIT distance="200" swimtime="00:01:47.80" />
                    <SPLIT distance="225" swimtime="00:01:58.32" />
                    <SPLIT distance="250" swimtime="00:02:11.06" />
                    <SPLIT distance="275" swimtime="00:02:24.39" />
                    <SPLIT distance="300" swimtime="00:02:38.12" />
                    <SPLIT distance="325" swimtime="00:02:48.36" />
                    <SPLIT distance="350" swimtime="00:03:00.43" />
                    <SPLIT distance="375" swimtime="00:03:12.90" />
                    <SPLIT distance="400" swimtime="00:03:25.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202663" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="163641" reactiontime="+39" />
                    <RELAYPOSITION number="3" athleteid="202666" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="120880" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Australia">
              <RESULTS>
                <RESULT eventid="132" place="2" lane="6" heat="1" swimtime="00:06:46.54" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:23.84" />
                    <SPLIT distance="75" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:00:49.33" />
                    <SPLIT distance="125" swimtime="00:01:02.26" />
                    <SPLIT distance="150" swimtime="00:01:15.37" />
                    <SPLIT distance="175" swimtime="00:01:28.65" />
                    <SPLIT distance="200" swimtime="00:01:41.50" />
                    <SPLIT distance="225" swimtime="00:01:52.18" />
                    <SPLIT distance="250" swimtime="00:02:04.53" />
                    <SPLIT distance="275" swimtime="00:02:17.17" />
                    <SPLIT distance="300" swimtime="00:02:30.03" />
                    <SPLIT distance="325" swimtime="00:02:42.85" />
                    <SPLIT distance="350" swimtime="00:02:56.06" />
                    <SPLIT distance="375" swimtime="00:03:09.10" />
                    <SPLIT distance="400" swimtime="00:03:21.85" />
                    <SPLIT distance="425" swimtime="00:03:32.38" />
                    <SPLIT distance="450" swimtime="00:03:45.11" />
                    <SPLIT distance="475" swimtime="00:03:58.16" />
                    <SPLIT distance="500" swimtime="00:04:11.15" />
                    <SPLIT distance="525" swimtime="00:04:24.04" />
                    <SPLIT distance="550" swimtime="00:04:37.42" />
                    <SPLIT distance="575" swimtime="00:04:50.48" />
                    <SPLIT distance="600" swimtime="00:05:03.35" />
                    <SPLIT distance="625" swimtime="00:05:14.23" />
                    <SPLIT distance="650" swimtime="00:05:27.05" />
                    <SPLIT distance="675" swimtime="00:05:40.08" />
                    <SPLIT distance="700" swimtime="00:05:53.18" />
                    <SPLIT distance="725" swimtime="00:06:06.40" />
                    <SPLIT distance="750" swimtime="00:06:19.93" />
                    <SPLIT distance="775" swimtime="00:06:33.41" />
                    <SPLIT distance="800" swimtime="00:06:46.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="163637" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="120880" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="202662" reactiontime="+6" />
                    <RELAYPOSITION number="4" athleteid="110896" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="4" lane="3" heat="2" swimtime="00:06:54.83" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.51" />
                    <SPLIT distance="50" swimtime="00:00:24.30" />
                    <SPLIT distance="75" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:00:50.50" />
                    <SPLIT distance="125" swimtime="00:01:03.88" />
                    <SPLIT distance="150" swimtime="00:01:17.26" />
                    <SPLIT distance="175" swimtime="00:01:30.88" />
                    <SPLIT distance="200" swimtime="00:01:44.33" />
                    <SPLIT distance="225" swimtime="00:01:55.06" />
                    <SPLIT distance="250" swimtime="00:02:07.62" />
                    <SPLIT distance="275" swimtime="00:02:20.74" />
                    <SPLIT distance="300" swimtime="00:02:33.71" />
                    <SPLIT distance="325" swimtime="00:02:46.80" />
                    <SPLIT distance="350" swimtime="00:03:00.31" />
                    <SPLIT distance="375" swimtime="00:03:13.71" />
                    <SPLIT distance="400" swimtime="00:03:26.53" />
                    <SPLIT distance="425" swimtime="00:03:37.60" />
                    <SPLIT distance="450" swimtime="00:03:50.31" />
                    <SPLIT distance="475" swimtime="00:04:03.40" />
                    <SPLIT distance="500" swimtime="00:04:16.70" />
                    <SPLIT distance="525" swimtime="00:04:30.13" />
                    <SPLIT distance="550" swimtime="00:04:43.62" />
                    <SPLIT distance="575" swimtime="00:04:57.32" />
                    <SPLIT distance="600" swimtime="00:05:10.90" />
                    <SPLIT distance="625" swimtime="00:05:22.17" />
                    <SPLIT distance="650" swimtime="00:05:34.97" />
                    <SPLIT distance="675" swimtime="00:05:48.07" />
                    <SPLIT distance="700" swimtime="00:06:01.36" />
                    <SPLIT distance="725" swimtime="00:06:14.73" />
                    <SPLIT distance="750" swimtime="00:06:28.16" />
                    <SPLIT distance="775" swimtime="00:06:41.91" />
                    <SPLIT distance="800" swimtime="00:06:54.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="120888" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="202662" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="150388" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="202654" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Australia">
              <RESULTS>
                <RESULT eventid="126" place="1" lane="2" heat="1" swimtime="00:01:23.44" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:21.25" />
                    <SPLIT distance="75" swimtime="00:00:30.98" />
                    <SPLIT distance="100" swimtime="00:00:42.00" />
                    <SPLIT distance="125" swimtime="00:00:52.09" />
                    <SPLIT distance="150" swimtime="00:01:03.10" />
                    <SPLIT distance="175" swimtime="00:01:12.69" />
                    <SPLIT distance="200" swimtime="00:01:23.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202663" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="156743" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="202662" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="120880" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="5" lane="1" heat="1" swimtime="00:01:24.42" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.34" />
                    <SPLIT distance="50" swimtime="00:00:21.24" />
                    <SPLIT distance="75" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:00:42.63" />
                    <SPLIT distance="125" swimtime="00:00:52.53" />
                    <SPLIT distance="150" swimtime="00:01:03.71" />
                    <SPLIT distance="175" swimtime="00:01:13.37" />
                    <SPLIT distance="200" swimtime="00:01:24.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202663" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="120878" reactiontime="+35" />
                    <RELAYPOSITION number="3" athleteid="202662" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="156743" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Australia">
              <RESULTS>
                <RESULT eventid="127" place="2" lane="5" heat="1" swimtime="00:01:28.03" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.07" />
                    <SPLIT distance="50" swimtime="00:00:20.97" />
                    <SPLIT distance="75" swimtime="00:00:30.65" />
                    <SPLIT distance="100" swimtime="00:00:41.68" />
                    <SPLIT distance="125" swimtime="00:00:53.10" />
                    <SPLIT distance="150" swimtime="00:01:05.41" />
                    <SPLIT distance="175" swimtime="00:01:16.13" />
                    <SPLIT distance="200" swimtime="00:01:28.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="120880" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="156743" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="173958" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="100650" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="2" lane="2" heat="1" swimtime="00:01:29.82" reactiontime="+71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.78" />
                    <SPLIT distance="50" swimtime="00:00:22.04" />
                    <SPLIT distance="75" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:00:43.01" />
                    <SPLIT distance="125" swimtime="00:00:54.41" />
                    <SPLIT distance="150" swimtime="00:01:06.84" />
                    <SPLIT distance="175" swimtime="00:01:17.70" />
                    <SPLIT distance="200" swimtime="00:01:29.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202662" reactiontime="+71" />
                    <RELAYPOSITION number="2" athleteid="156743" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="105256" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="100650" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Australia">
              <RESULTS>
                <RESULT eventid="108" place="1" lane="4" heat="1" swimtime="00:03:25.43" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:25.28" />
                    <SPLIT distance="75" swimtime="00:00:38.79" />
                    <SPLIT distance="100" swimtime="00:00:52.19" />
                    <SPLIT distance="125" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:16.83" />
                    <SPLIT distance="175" swimtime="00:01:30.18" />
                    <SPLIT distance="200" swimtime="00:01:43.47" />
                    <SPLIT distance="225" swimtime="00:01:55.04" />
                    <SPLIT distance="250" swimtime="00:02:08.34" />
                    <SPLIT distance="275" swimtime="00:02:21.91" />
                    <SPLIT distance="300" swimtime="00:02:35.47" />
                    <SPLIT distance="325" swimtime="00:02:46.59" />
                    <SPLIT distance="350" swimtime="00:02:59.36" />
                    <SPLIT distance="375" swimtime="00:03:12.47" />
                    <SPLIT distance="400" swimtime="00:03:25.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="163620" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="105256" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="173958" reactiontime="+45" />
                    <RELAYPOSITION number="4" athleteid="100650" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="1" lane="3" heat="2" swimtime="00:03:28.58" reactiontime="+71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:25.06" />
                    <SPLIT distance="75" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:00:52.11" />
                    <SPLIT distance="125" swimtime="00:01:03.66" />
                    <SPLIT distance="150" swimtime="00:01:17.03" />
                    <SPLIT distance="175" swimtime="00:01:30.35" />
                    <SPLIT distance="200" swimtime="00:01:43.54" />
                    <SPLIT distance="225" swimtime="00:01:55.68" />
                    <SPLIT distance="250" swimtime="00:02:09.27" />
                    <SPLIT distance="275" swimtime="00:02:23.30" />
                    <SPLIT distance="300" swimtime="00:02:36.82" />
                    <SPLIT distance="325" swimtime="00:02:48.24" />
                    <SPLIT distance="350" swimtime="00:03:01.35" />
                    <SPLIT distance="375" swimtime="00:03:14.98" />
                    <SPLIT distance="400" swimtime="00:03:28.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="173958" reactiontime="+71" />
                    <RELAYPOSITION number="2" athleteid="105256" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="111247" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="100650" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Australia">
              <RESULTS>
                <RESULT eventid="147" place="2" lane="5" heat="1" swimtime="00:03:44.92" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="75" swimtime="00:00:41.40" />
                    <SPLIT distance="100" swimtime="00:00:55.74" />
                    <SPLIT distance="125" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:25.59" />
                    <SPLIT distance="175" swimtime="00:01:42.58" />
                    <SPLIT distance="200" swimtime="00:02:00.23" />
                    <SPLIT distance="225" swimtime="00:02:11.41" />
                    <SPLIT distance="250" swimtime="00:02:25.11" />
                    <SPLIT distance="275" swimtime="00:02:39.31" />
                    <SPLIT distance="300" swimtime="00:02:54.16" />
                    <SPLIT distance="325" swimtime="00:03:05.41" />
                    <SPLIT distance="350" swimtime="00:03:18.30" />
                    <SPLIT distance="375" swimtime="00:03:31.76" />
                    <SPLIT distance="400" swimtime="00:03:44.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130172" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="129244" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="100650" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="173958" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="2" lane="3" heat="1" swimtime="00:03:48.90" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                    <SPLIT distance="75" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:00:55.81" />
                    <SPLIT distance="125" swimtime="00:01:09.35" />
                    <SPLIT distance="150" swimtime="00:01:25.99" />
                    <SPLIT distance="175" swimtime="00:01:43.34" />
                    <SPLIT distance="200" swimtime="00:02:01.05" />
                    <SPLIT distance="225" swimtime="00:02:12.67" />
                    <SPLIT distance="250" swimtime="00:02:27.05" />
                    <SPLIT distance="275" swimtime="00:02:41.85" />
                    <SPLIT distance="300" swimtime="00:02:57.32" />
                    <SPLIT distance="325" swimtime="00:03:08.95" />
                    <SPLIT distance="350" swimtime="00:03:22.11" />
                    <SPLIT distance="375" swimtime="00:03:35.51" />
                    <SPLIT distance="400" swimtime="00:03:48.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="163620" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="150358" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="202753" reactiontime="+22" />
                    <RELAYPOSITION number="4" athleteid="173958" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Australia">
              <RESULTS>
                <RESULT eventid="117" place="1" lane="5" heat="1" swimtime="00:07:30.87" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:26.50" />
                    <SPLIT distance="75" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:00:55.10" />
                    <SPLIT distance="125" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:24.17" />
                    <SPLIT distance="175" swimtime="00:01:38.70" />
                    <SPLIT distance="200" swimtime="00:01:53.13" />
                    <SPLIT distance="225" swimtime="00:02:05.62" />
                    <SPLIT distance="250" swimtime="00:02:19.66" />
                    <SPLIT distance="275" swimtime="00:02:34.07" />
                    <SPLIT distance="300" swimtime="00:02:48.57" />
                    <SPLIT distance="325" swimtime="00:03:02.98" />
                    <SPLIT distance="350" swimtime="00:03:17.60" />
                    <SPLIT distance="375" swimtime="00:03:32.09" />
                    <SPLIT distance="400" swimtime="00:03:45.96" />
                    <SPLIT distance="425" swimtime="00:03:58.13" />
                    <SPLIT distance="450" swimtime="00:04:12.09" />
                    <SPLIT distance="475" swimtime="00:04:26.28" />
                    <SPLIT distance="500" swimtime="00:04:40.60" />
                    <SPLIT distance="525" swimtime="00:04:55.01" />
                    <SPLIT distance="550" swimtime="00:05:09.51" />
                    <SPLIT distance="575" swimtime="00:05:24.22" />
                    <SPLIT distance="600" swimtime="00:05:38.63" />
                    <SPLIT distance="625" swimtime="00:05:50.64" />
                    <SPLIT distance="650" swimtime="00:06:04.52" />
                    <SPLIT distance="675" swimtime="00:06:18.74" />
                    <SPLIT distance="700" swimtime="00:06:32.96" />
                    <SPLIT distance="725" swimtime="00:06:47.40" />
                    <SPLIT distance="750" swimtime="00:07:01.94" />
                    <SPLIT distance="775" swimtime="00:07:16.58" />
                    <SPLIT distance="800" swimtime="00:07:30.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="105256" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="163620" reactiontime="+41" />
                    <RELAYPOSITION number="3" athleteid="111247" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="150371" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="2" lane="5" heat="2" swimtime="00:07:44.77" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.74" />
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="75" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:00:56.53" />
                    <SPLIT distance="125" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:26.27" />
                    <SPLIT distance="175" swimtime="00:01:41.39" />
                    <SPLIT distance="200" swimtime="00:01:55.85" />
                    <SPLIT distance="225" swimtime="00:02:08.10" />
                    <SPLIT distance="250" swimtime="00:02:22.15" />
                    <SPLIT distance="275" swimtime="00:02:36.65" />
                    <SPLIT distance="300" swimtime="00:02:51.41" />
                    <SPLIT distance="325" swimtime="00:03:05.99" />
                    <SPLIT distance="350" swimtime="00:03:20.74" />
                    <SPLIT distance="375" swimtime="00:03:35.62" />
                    <SPLIT distance="400" swimtime="00:03:50.11" />
                    <SPLIT distance="425" swimtime="00:04:02.84" />
                    <SPLIT distance="450" swimtime="00:04:17.52" />
                    <SPLIT distance="475" swimtime="00:04:32.33" />
                    <SPLIT distance="500" swimtime="00:04:47.10" />
                    <SPLIT distance="525" swimtime="00:05:01.93" />
                    <SPLIT distance="550" swimtime="00:05:16.91" />
                    <SPLIT distance="575" swimtime="00:05:31.83" />
                    <SPLIT distance="600" swimtime="00:05:46.28" />
                    <SPLIT distance="625" swimtime="00:05:59.06" />
                    <SPLIT distance="650" swimtime="00:06:13.65" />
                    <SPLIT distance="675" swimtime="00:06:28.60" />
                    <SPLIT distance="700" swimtime="00:06:43.80" />
                    <SPLIT distance="725" swimtime="00:06:59.27" />
                    <SPLIT distance="750" swimtime="00:07:14.53" />
                    <SPLIT distance="775" swimtime="00:07:29.92" />
                    <SPLIT distance="800" swimtime="00:07:44.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="111247" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="173958" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="172303" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="161731" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Australia">
              <RESULTS>
                <RESULT eventid="125" place="2" lane="5" heat="1" swimtime="00:01:34.23" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.77" />
                    <SPLIT distance="50" swimtime="00:00:23.98" />
                    <SPLIT distance="75" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:00:47.49" />
                    <SPLIT distance="125" swimtime="00:00:59.12" />
                    <SPLIT distance="150" swimtime="00:01:11.50" />
                    <SPLIT distance="175" swimtime="00:01:22.34" />
                    <SPLIT distance="200" swimtime="00:01:34.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="173958" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="105256" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="163620" reactiontime="+52" />
                    <RELAYPOSITION number="4" athleteid="100650" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="2" lane="6" heat="1" swimtime="00:01:36.14" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:23.85" />
                    <SPLIT distance="75" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:00:47.95" />
                    <SPLIT distance="125" swimtime="00:00:59.51" />
                    <SPLIT distance="150" swimtime="00:01:12.24" />
                    <SPLIT distance="175" swimtime="00:01:23.81" />
                    <SPLIT distance="200" swimtime="00:01:36.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="173958" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="202753" reactiontime="+30" />
                    <RELAYPOSITION number="3" athleteid="172303" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="163620" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Australia">
              <RESULTS>
                <RESULT eventid="134" place="1" lane="4" heat="1" swimtime="00:01:42.35" reactiontime="+52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                    <SPLIT distance="50" swimtime="00:00:25.49" />
                    <SPLIT distance="75" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:00:54.60" />
                    <SPLIT distance="125" swimtime="00:01:05.57" />
                    <SPLIT distance="150" swimtime="00:01:19.03" />
                    <SPLIT distance="175" swimtime="00:01:30.21" />
                    <SPLIT distance="200" swimtime="00:01:42.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="163620" reactiontime="+52" />
                    <RELAYPOSITION number="2" athleteid="150358" reactiontime="+27" />
                    <RELAYPOSITION number="3" athleteid="100650" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="105256" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="1" lane="8" heat="1" swimtime="00:01:44.78" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                    <SPLIT distance="75" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:00:56.63" />
                    <SPLIT distance="125" swimtime="00:01:07.73" />
                    <SPLIT distance="150" swimtime="00:01:21.42" />
                    <SPLIT distance="175" swimtime="00:01:32.63" />
                    <SPLIT distance="200" swimtime="00:01:44.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130172" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="129244" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="100650" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="105256" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Australia">
              <RESULTS>
                <RESULT eventid="11" place="10" lane="8" heat="1" swimtime="00:01:39.41" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:23.87" />
                    <SPLIT distance="75" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:00:50.04" />
                    <SPLIT distance="125" swimtime="00:01:01.48" />
                    <SPLIT distance="150" swimtime="00:01:15.55" />
                    <SPLIT distance="175" swimtime="00:01:27.03" />
                    <SPLIT distance="200" swimtime="00:01:39.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="120897" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="120878" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="202753" reactiontime="+21" />
                    <RELAYPOSITION number="4" athleteid="173958" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Australia">
              <RESULTS>
                <RESULT eventid="135" place="3" lane="1" heat="1" swimtime="00:01:30.81" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.04" />
                    <SPLIT distance="50" swimtime="00:00:22.66" />
                    <SPLIT distance="75" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:00:48.58" />
                    <SPLIT distance="125" swimtime="00:00:58.39" />
                    <SPLIT distance="150" swimtime="00:01:10.33" />
                    <SPLIT distance="175" swimtime="00:01:20.06" />
                    <SPLIT distance="200" swimtime="00:01:30.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202663" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="120878" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="156743" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="120880" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="7" lane="6" heat="2" swimtime="00:01:33.25" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:22.95" />
                    <SPLIT distance="75" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:00:49.25" />
                    <SPLIT distance="125" swimtime="00:00:59.56" />
                    <SPLIT distance="150" swimtime="00:01:11.97" />
                    <SPLIT distance="175" swimtime="00:01:22.06" />
                    <SPLIT distance="200" swimtime="00:01:33.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202663" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="120878" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="202666" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="202662" reactiontime="+6" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Austria" shortname="AUT" code="AUT" nation="AUT" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="106854" lastname="REITSHAMMER" firstname="Bernhard" gender="M" birthdate="1994-06-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.80" eventid="16" heat="7" lane="3">
                  <MEETINFO date="2021-11-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.10" eventid="41" heat="8" lane="3">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.91" eventid="23" heat="4" lane="3">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="11" lane="3" heat="7" heatid="70016" swimtime="00:00:57.66" reactiontime="+68" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                    <SPLIT distance="75" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:00:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="15" lane="7" heat="2" heatid="20216" swimtime="00:00:57.98" reactiontime="+66" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                    <SPLIT distance="75" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:00:57.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="18" lane="3" heat="8" heatid="80041" swimtime="00:00:26.64" reactiontime="+67" points="821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="7" lane="1" heat="1" heatid="10123" swimtime="00:00:52.01" reactiontime="+66" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.77" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                    <SPLIT distance="75" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:00:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="8" lane="3" heat="4" heatid="40023" swimtime="00:00:52.28" reactiontime="+67" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.84" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                    <SPLIT distance="75" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:00:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="7" lane="6" heat="1" heatid="10223" swimtime="00:00:51.78" reactiontime="+67" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.85" />
                    <SPLIT distance="50" swimtime="00:00:23.85" />
                    <SPLIT distance="75" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:00:51.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154837" lastname="BUCHER" firstname="Simon" gender="M" birthdate="2000-05-23">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.70" eventid="39" heat="8" lane="6">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.58" eventid="19" heat="5" lane="7">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.70" eventid="5" heat="9" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="6" lane="7" heat="1" heatid="10139" swimtime="00:00:49.39" reactiontime="+59" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.41" />
                    <SPLIT distance="50" swimtime="00:00:23.08" />
                    <SPLIT distance="75" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:00:49.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="8" lane="6" heat="8" heatid="80039" swimtime="00:00:50.06" reactiontime="+61" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.52" />
                    <SPLIT distance="50" swimtime="00:00:23.27" />
                    <SPLIT distance="75" swimtime="00:00:36.62" />
                    <SPLIT distance="100" swimtime="00:00:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="6" lane="6" heat="1" heatid="10239" swimtime="00:00:49.72" reactiontime="+59" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.46" />
                    <SPLIT distance="50" swimtime="00:00:23.08" />
                    <SPLIT distance="75" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:00:49.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="19" lane="7" heat="5" heatid="50019" swimtime="00:00:23.55" reactiontime="+57" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:23.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="13" lane="1" heat="9" heatid="90005" swimtime="00:00:22.44" reactiontime="+59" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:22.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="11" lane="1" heat="2" heatid="20205" swimtime="00:00:22.35" reactiontime="+61" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.29" />
                    <SPLIT distance="50" swimtime="00:00:22.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149509" lastname="GIGLER" firstname="Heiko" gender="M" birthdate="1996-06-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.74" eventid="14" heat="10" lane="6">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.25" eventid="31" heat="11" lane="7">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.04" eventid="23" heat="5" lane="6">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="10" lane="6" heat="10" heatid="100014" swimtime="00:00:46.64" reactiontime="+62" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:22.16" />
                    <SPLIT distance="75" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:00:46.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="14" lane="2" heat="1" heatid="10214" swimtime="00:00:46.92" reactiontime="+62" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.46" />
                    <SPLIT distance="50" swimtime="00:00:22.14" />
                    <SPLIT distance="75" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:00:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="25" lane="7" heat="11" heatid="110031" swimtime="00:00:21.42" reactiontime="+62" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.33" />
                    <SPLIT distance="50" swimtime="00:00:21.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="12" lane="6" heat="5" heatid="50023" swimtime="00:00:52.58" reactiontime="+64" points="823">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.81" />
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                    <SPLIT distance="75" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:00:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="10" lane="1" heat="2" heatid="20223" swimtime="00:00:52.10" reactiontime="+63" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.64" />
                    <SPLIT distance="50" swimtime="00:00:23.45" />
                    <SPLIT distance="75" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:00:52.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="192888" lastname="HERCOG" firstname="Jan" gender="M" birthdate="1998-02-10">
              <ENTRIES>
                <ENTRY entrytime="00:14:56.68" eventid="10" heat="1" lane="4">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="15" lane="4" heat="1" heatid="10010" swimtime="00:15:00.36" reactiontime="+67" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                    <SPLIT distance="75" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:00:55.81" />
                    <SPLIT distance="125" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:25.16" />
                    <SPLIT distance="175" swimtime="00:01:39.91" />
                    <SPLIT distance="200" swimtime="00:01:54.55" />
                    <SPLIT distance="225" swimtime="00:02:09.34" />
                    <SPLIT distance="250" swimtime="00:02:24.22" />
                    <SPLIT distance="275" swimtime="00:02:39.05" />
                    <SPLIT distance="300" swimtime="00:02:53.97" />
                    <SPLIT distance="325" swimtime="00:03:08.68" />
                    <SPLIT distance="350" swimtime="00:03:23.51" />
                    <SPLIT distance="375" swimtime="00:03:38.34" />
                    <SPLIT distance="400" swimtime="00:03:53.32" />
                    <SPLIT distance="425" swimtime="00:04:08.16" />
                    <SPLIT distance="450" swimtime="00:04:23.17" />
                    <SPLIT distance="475" swimtime="00:04:38.06" />
                    <SPLIT distance="500" swimtime="00:04:53.04" />
                    <SPLIT distance="525" swimtime="00:05:07.97" />
                    <SPLIT distance="550" swimtime="00:05:22.90" />
                    <SPLIT distance="575" swimtime="00:05:37.98" />
                    <SPLIT distance="600" swimtime="00:05:52.92" />
                    <SPLIT distance="625" swimtime="00:06:07.92" />
                    <SPLIT distance="650" swimtime="00:06:23.00" />
                    <SPLIT distance="675" swimtime="00:06:38.13" />
                    <SPLIT distance="700" swimtime="00:06:53.21" />
                    <SPLIT distance="725" swimtime="00:07:08.51" />
                    <SPLIT distance="750" swimtime="00:07:23.60" />
                    <SPLIT distance="775" swimtime="00:07:38.90" />
                    <SPLIT distance="800" swimtime="00:07:53.96" />
                    <SPLIT distance="825" swimtime="00:08:09.16" />
                    <SPLIT distance="850" swimtime="00:08:24.22" />
                    <SPLIT distance="875" swimtime="00:08:39.43" />
                    <SPLIT distance="900" swimtime="00:08:54.56" />
                    <SPLIT distance="925" swimtime="00:09:09.82" />
                    <SPLIT distance="950" swimtime="00:09:24.95" />
                    <SPLIT distance="975" swimtime="00:09:40.24" />
                    <SPLIT distance="1000" swimtime="00:09:55.51" />
                    <SPLIT distance="1025" swimtime="00:10:10.89" />
                    <SPLIT distance="1050" swimtime="00:10:26.05" />
                    <SPLIT distance="1075" swimtime="00:10:41.37" />
                    <SPLIT distance="1100" swimtime="00:10:56.56" />
                    <SPLIT distance="1125" swimtime="00:11:11.85" />
                    <SPLIT distance="1150" swimtime="00:11:27.06" />
                    <SPLIT distance="1175" swimtime="00:11:42.41" />
                    <SPLIT distance="1200" swimtime="00:11:57.58" />
                    <SPLIT distance="1225" swimtime="00:12:12.84" />
                    <SPLIT distance="1250" swimtime="00:12:28.00" />
                    <SPLIT distance="1275" swimtime="00:12:43.21" />
                    <SPLIT distance="1300" swimtime="00:12:58.36" />
                    <SPLIT distance="1325" swimtime="00:13:13.62" />
                    <SPLIT distance="1350" swimtime="00:13:28.94" />
                    <SPLIT distance="1375" swimtime="00:13:44.26" />
                    <SPLIT distance="1400" swimtime="00:13:59.50" />
                    <SPLIT distance="1425" swimtime="00:14:14.82" />
                    <SPLIT distance="1450" swimtime="00:14:30.23" />
                    <SPLIT distance="1475" swimtime="00:14:45.57" />
                    <SPLIT distance="1500" swimtime="00:15:00.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125412" lastname="PILHATSCH" firstname="Caroline" gender="F" birthdate="1999-03-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.43" eventid="2" heat="4" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.05" eventid="18" heat="7" lane="3">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="29" lane="1" heat="4" heatid="40002" swimtime="00:00:59.71" reactiontime="+59" points="776">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:00:59.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="21" lane="3" heat="7" heatid="70018" swimtime="00:00:26.81" reactiontime="+56" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105517" lastname="KREUNDL" firstname="Lena" gender="F" birthdate="1997-09-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.82" eventid="15" heat="4" lane="3">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.39" eventid="13" heat="8" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.51" eventid="28" heat="2" lane="4">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.76" eventid="6" heat="3" lane="7">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.08" eventid="22" heat="2" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="32" lane="3" heat="4" heatid="40015" swimtime="00:01:07.15" reactiontime="+68" points="800">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.44" />
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="75" swimtime="00:00:49.15" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="20" lane="1" heat="8" heatid="80013" swimtime="00:00:53.67" reactiontime="+65" points="820">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="75" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:00:53.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="-1" lane="4" heat="2" heatid="20028" swimtime="NT" status="DNS" />
                <RESULT eventid="6" place="14" lane="7" heat="3" heatid="30006" swimtime="00:02:08.44" reactiontime="+68" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="75" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:00.30" />
                    <SPLIT distance="125" swimtime="00:01:18.64" />
                    <SPLIT distance="150" swimtime="00:01:37.23" />
                    <SPLIT distance="175" swimtime="00:01:53.34" />
                    <SPLIT distance="200" swimtime="00:02:08.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="7" lane="7" heat="1" heatid="10122" swimtime="00:00:58.79" reactiontime="+66" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                    <SPLIT distance="75" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:00:58.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="7" lane="3" heat="2" heatid="20022" swimtime="00:00:59.29" reactiontime="+67" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="75" swimtime="00:00:44.80" />
                    <SPLIT distance="100" swimtime="00:00:59.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="6" lane="6" heat="2" heatid="20222" swimtime="00:00:59.04" reactiontime="+65" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                    <SPLIT distance="75" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:00:59.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Austria">
              <RESULTS>
                <RESULT eventid="11" place="12" lane="5" heat="2" swimtime="00:01:39.71" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.21" />
                    <SPLIT distance="50" swimtime="00:00:27.06" />
                    <SPLIT distance="75" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:00:52.85" />
                    <SPLIT distance="125" swimtime="00:01:02.83" />
                    <SPLIT distance="150" swimtime="00:01:15.19" />
                    <SPLIT distance="175" swimtime="00:01:26.79" />
                    <SPLIT distance="200" swimtime="00:01:39.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="125412" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="106854" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="154837" reactiontime="+15" />
                    <RELAYPOSITION number="4" athleteid="105517" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Bahamas" shortname="BAH" code="BAH" nation="BAH" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="162306" lastname="TAYLOR" firstname="Lamar" gender="M" birthdate="2003-06-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.25" eventid="14" heat="5" lane="4">
                  <MEETINFO date="2022-07-09" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.38" eventid="19" heat="3" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.21" eventid="5" heat="4" lane="3">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.45" eventid="31" heat="6" lane="2">
                  <MEETINFO date="2022-08-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="36" lane="4" heat="5" heatid="50014" swimtime="00:00:47.76" reactiontime="+60" points="827">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.49" />
                    <SPLIT distance="75" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:00:47.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="20" lane="3" heat="3" heatid="30019" swimtime="00:00:23.58" reactiontime="+59" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                    <SPLIT distance="50" swimtime="00:00:23.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="-1" lane="3" heat="4" heatid="40005" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="28" lane="2" heat="6" heatid="60031" swimtime="00:00:21.45" reactiontime="+61" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.38" />
                    <SPLIT distance="50" swimtime="00:00:21.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213102" lastname="THOMPSON" firstname="Luke Kennedy" gender="M" birthdate="2001-08-03">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.44" eventid="44" heat="1" lane="5">
                  <MEETINFO date="2022-07-30" />
                </ENTRY>
                <ENTRY entrytime="00:04:04.90" eventid="24" heat="1" lane="6">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="40" lane="5" heat="1" heatid="10044" swimtime="00:01:51.31" reactiontime="+60" points="711">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="75" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="125" swimtime="00:01:08.88" />
                    <SPLIT distance="150" swimtime="00:01:23.16" />
                    <SPLIT distance="175" swimtime="00:01:37.70" />
                    <SPLIT distance="200" swimtime="00:01:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="28" lane="6" heat="1" heatid="10024" swimtime="00:03:56.22" reactiontime="+60" points="725">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                    <SPLIT distance="50" swimtime="00:00:26.70" />
                    <SPLIT distance="75" swimtime="00:00:41.17" />
                    <SPLIT distance="100" swimtime="00:00:55.90" />
                    <SPLIT distance="125" swimtime="00:01:10.73" />
                    <SPLIT distance="150" swimtime="00:01:25.48" />
                    <SPLIT distance="175" swimtime="00:01:40.44" />
                    <SPLIT distance="200" swimtime="00:01:55.66" />
                    <SPLIT distance="225" swimtime="00:02:10.64" />
                    <SPLIT distance="250" swimtime="00:02:25.87" />
                    <SPLIT distance="275" swimtime="00:02:40.80" />
                    <SPLIT distance="300" swimtime="00:02:56.02" />
                    <SPLIT distance="325" swimtime="00:03:11.24" />
                    <SPLIT distance="350" swimtime="00:03:26.47" />
                    <SPLIT distance="375" swimtime="00:03:41.91" />
                    <SPLIT distance="400" swimtime="00:03:56.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108581" lastname="RUSSELL" firstname="Victoria" gender="F" birthdate="2000-07-26">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:14.97" eventid="15" heat="2" lane="5">
                  <MEETINFO date="2022-04-10" />
                </ENTRY>
                <ENTRY entrytime="00:00:33.68" eventid="40" heat="3" lane="3">
                  <MEETINFO date="2022-07-09" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="40" lane="5" heat="2" heatid="20015" swimtime="00:01:11.56" reactiontime="+75" points="661">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.46" />
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="75" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="30" lane="3" heat="3" heatid="30040" swimtime="00:00:32.54" reactiontime="+70" points="676">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.91" />
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="203180" lastname="GIBBS" firstname="Rhaniska" gender="F" birthdate="2006-04-19">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:28.62" eventid="4" heat="3" lane="7">
                  <MEETINFO date="2022-07-08" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.68" eventid="30" heat="4" lane="7">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="31" lane="7" heat="3" heatid="30004" swimtime="00:00:28.07" reactiontime="+61" points="655">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="35" lane="7" heat="4" heatid="40030" swimtime="00:00:26.16" reactiontime="+61" points="673">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Bahamas">
              <RESULTS>
                <RESULT eventid="27" place="16" lane="6" heat="4" swimtime="00:01:36.95" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:21.65" />
                    <SPLIT distance="75" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:00:44.95" />
                    <SPLIT distance="125" swimtime="00:00:57.00" />
                    <SPLIT distance="150" swimtime="00:01:10.65" />
                    <SPLIT distance="175" swimtime="00:01:23.32" />
                    <SPLIT distance="200" swimtime="00:01:36.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="162306" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="213102" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="203180" reactiontime="-3" />
                    <RELAYPOSITION number="4" athleteid="108581" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Bahamas">
              <RESULTS>
                <RESULT eventid="11" place="22" lane="7" heat="3" swimtime="00:01:46.93" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:24.19" />
                    <SPLIT distance="75" swimtime="00:00:38.79" />
                    <SPLIT distance="100" swimtime="00:00:56.47" />
                    <SPLIT distance="125" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:20.97" />
                    <SPLIT distance="175" swimtime="00:01:33.50" />
                    <SPLIT distance="200" swimtime="00:01:46.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="162306" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="108581" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="213102" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="203180" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Bangladesh" shortname="BAN" code="BAN" nation="BAN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197102" lastname="REZA" firstname="Md Asif" gender="M" birthdate="1996-10-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.24" eventid="14" heat="3" lane="1">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.28" eventid="31" heat="4" lane="4">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="67" lane="1" heat="3" heatid="30014" swimtime="00:00:52.91" reactiontime="+64" points="608">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.06" />
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                    <SPLIT distance="75" swimtime="00:00:39.16" />
                    <SPLIT distance="100" swimtime="00:00:52.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="59" lane="4" heat="4" heatid="40031" swimtime="00:00:24.24" reactiontime="+68" points="575">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.81" />
                    <SPLIT distance="50" swimtime="00:00:24.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105108" lastname="AKTAR" firstname="Sonia" gender="F" birthdate="1997-07-15">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="13" heat="1" lane="5" />
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="59" lane="5" heat="1" heatid="10013" swimtime="00:01:05.05" reactiontime="+70" points="460">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="75" swimtime="00:00:48.58" />
                    <SPLIT distance="100" swimtime="00:01:05.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="50" lane="7" heat="1" heatid="10030" swimtime="00:00:29.75" reactiontime="+72" points="457">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.75" />
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Barbados" shortname="BAR" code="BAR" nation="BAR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="211014" lastname="CHEE-A-TOW" firstname="Jake" gender="M" birthdate="2004-10-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.37" eventid="14" heat="2" lane="4">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.34" eventid="21" heat="1" lane="4">
                  <MEETINFO date="2022-07-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="72" lane="4" heat="2" heatid="20014" swimtime="00:00:53.62" reactiontime="+57" points="584">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                    <SPLIT distance="75" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:00:53.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="25" lane="4" heat="1" heatid="10021" swimtime="00:02:07.92" reactiontime="+57" points="605">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="75" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:00:59.43" />
                    <SPLIT distance="125" swimtime="00:01:16.13" />
                    <SPLIT distance="150" swimtime="00:01:33.06" />
                    <SPLIT distance="175" swimtime="00:01:50.43" />
                    <SPLIT distance="200" swimtime="00:02:07.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Burundi" shortname="BDI" code="BDI" nation="BDI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="130536" lastname="IRAKOZE" firstname="Carel Van Melvin" gender="M" birthdate="2000-10-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.39" eventid="3" heat="1" lane="4">
                  <MEETINFO date="2021-10-15" />
                </ENTRY>
                <ENTRY entrytime="00:01:14.88" eventid="16" heat="1" lane="6">
                  <MEETINFO date="2021-10-11" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="39" lane="4" heat="1" heatid="10003" swimtime="00:01:02.86" reactiontime="+70" points="454">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="75" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="59" lane="6" heat="1" heatid="10016" swimtime="00:01:10.11" reactiontime="+74" points="490">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.75" />
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="75" swimtime="00:00:50.03" />
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Belgium" shortname="BEL" code="BEL" nation="BEL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198045" lastname="GASPARD" firstname="Florine" gender="F" birthdate="2001-12-28">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.45" eventid="15" heat="7" lane="8">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.70" eventid="40" heat="7" lane="6">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="19" lane="8" heat="7" heatid="70015" swimtime="00:01:05.49" reactiontime="+66" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.92" />
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="75" swimtime="00:00:47.63" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="9" lane="6" heat="7" heatid="70040" swimtime="00:00:29.79" reactiontime="+66" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="11" lane="2" heat="2" heatid="20240" swimtime="00:00:29.98" reactiontime="+65" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165101" lastname="DUMONT" firstname="Valentine" gender="F" birthdate="2000-07-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.81" eventid="13" heat="8" lane="8">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.34" eventid="43" heat="4" lane="2">
                  <MEETINFO date="2021-11-21" />
                </ENTRY>
                <ENTRY entrytime="00:04:01.84" eventid="1" heat="4" lane="6">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="21" lane="8" heat="8" heatid="80013" swimtime="00:00:53.77" reactiontime="+70" points="816">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                    <SPLIT distance="75" swimtime="00:00:39.96" />
                    <SPLIT distance="100" swimtime="00:00:53.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="13" lane="2" heat="4" heatid="40043" swimtime="00:01:55.80" reactiontime="+71" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                    <SPLIT distance="75" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:00:56.00" />
                    <SPLIT distance="125" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:25.76" />
                    <SPLIT distance="175" swimtime="00:01:40.94" />
                    <SPLIT distance="200" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="12" lane="6" heat="4" heatid="40001" swimtime="00:04:07.37" reactiontime="+73" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="75" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:00:58.41" />
                    <SPLIT distance="125" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:01:28.97" />
                    <SPLIT distance="175" swimtime="00:01:44.44" />
                    <SPLIT distance="200" swimtime="00:02:00.07" />
                    <SPLIT distance="225" swimtime="00:02:15.86" />
                    <SPLIT distance="250" swimtime="00:02:31.62" />
                    <SPLIT distance="275" swimtime="00:02:47.38" />
                    <SPLIT distance="300" swimtime="00:03:03.34" />
                    <SPLIT distance="325" swimtime="00:03:19.40" />
                    <SPLIT distance="350" swimtime="00:03:35.71" />
                    <SPLIT distance="375" swimtime="00:03:51.96" />
                    <SPLIT distance="400" swimtime="00:04:07.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165204" lastname="VERMEIREN" firstname="Fleur" gender="F" birthdate="2002-06-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.22" eventid="40" heat="6" lane="1">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="15" lane="1" heat="6" heatid="60040" swimtime="00:00:30.22" reactiontime="+67" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.89" />
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="16" lane="8" heat="2" heatid="20240" swimtime="00:00:30.29" reactiontime="+69" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Benin" shortname="BEN" code="BEN" nation="BEN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197396" lastname="DANSOU" firstname="Marc Pascal Pierre" gender="M" birthdate="1983-11-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.06" eventid="14" heat="3" lane="3">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.06" eventid="41" heat="2" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="70" lane="3" heat="3" heatid="30014" swimtime="00:00:53.46" reactiontime="+64" points="590">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:25.31" />
                    <SPLIT distance="75" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:00:53.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="-1" lane="5" heat="2" heatid="20041" swimtime="00:00:29.50" status="DSQ" reactiontime="+65" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Bhutan" shortname="BHU" code="BHU" nation="BHU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="160613" lastname="LHENDUP" firstname="Kinley" gender="M" birthdate="2004-06-16">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="39" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="7" heat="1" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="52" lane="3" heat="1" heatid="10039" swimtime="00:01:00.99" reactiontime="+68" points="480">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="75" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:00.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="37" lane="2" heat="1" heatid="10007" swimtime="00:02:20.63" reactiontime="+68" points="473">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                    <SPLIT distance="75" swimtime="00:00:46.48" />
                    <SPLIT distance="100" swimtime="00:01:03.91" />
                    <SPLIT distance="125" swimtime="00:01:25.16" />
                    <SPLIT distance="150" swimtime="00:01:46.64" />
                    <SPLIT distance="175" swimtime="00:02:04.26" />
                    <SPLIT distance="200" swimtime="00:02:20.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160828" lastname="TENZIN" firstname="Sangay" gender="M" birthdate="2003-09-07">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="14" heat="1" lane="8" />
                <ENTRY entrytime="NT" eventid="44" heat="1" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="77" lane="8" heat="1" heatid="10014" swimtime="00:00:55.46" reactiontime="+65" points="528">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.50" />
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                    <SPLIT distance="75" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:00:55.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="45" lane="7" heat="1" heatid="10044" swimtime="00:02:03.80" reactiontime="+72" points="517">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="75" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:00:59.85" />
                    <SPLIT distance="125" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:31.95" />
                    <SPLIT distance="175" swimtime="00:01:48.07" />
                    <SPLIT distance="200" swimtime="00:02:03.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Bosnia Herzegovina" shortname="BIH" code="BIH" nation="BIH" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="117160" lastname="MESETOVIC" firstname="Adi" gender="M" birthdate="1997-04-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.46" eventid="14" heat="5" lane="6">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.78" eventid="31" heat="5" lane="4">
                  <MEETINFO date="2022-08-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="46" lane="6" heat="5" heatid="50014" swimtime="00:00:48.97" reactiontime="+66" points="767">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.94" />
                    <SPLIT distance="50" swimtime="00:00:23.34" />
                    <SPLIT distance="75" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:00:48.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="46" lane="4" heat="5" heatid="50031" swimtime="00:00:22.27" reactiontime="+65" points="741">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197064" lastname="PUDAR" firstname="Lana" gender="F" birthdate="2006-01-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.28" eventid="38" heat="2" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.05" eventid="13" heat="6" lane="2">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.88" eventid="20" heat="3" lane="5">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="9" lane="5" heat="2" heatid="20038" swimtime="00:00:56.89" reactiontime="+71" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.25" />
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                    <SPLIT distance="75" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:00:56.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="10" lane="2" heat="2" heatid="20238" swimtime="00:00:56.71" reactiontime="+70" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="75" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:00:56.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="33" lane="2" heat="6" heatid="60013" swimtime="00:00:54.76" reactiontime="+68" points="772">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.72" />
                    <SPLIT distance="50" swimtime="00:00:26.63" />
                    <SPLIT distance="75" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:00:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="120" place="5" lane="8" heat="1" heatid="10120" swimtime="00:02:05.23" reactiontime="+74" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.66" />
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="75" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:00:59.97" />
                    <SPLIT distance="125" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:32.51" />
                    <SPLIT distance="175" swimtime="00:01:48.78" />
                    <SPLIT distance="200" swimtime="00:02:05.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="8" lane="5" heat="3" heatid="30020" swimtime="00:02:05.87" reactiontime="+74" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="75" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="125" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:32.77" />
                    <SPLIT distance="175" swimtime="00:01:49.18" />
                    <SPLIT distance="200" swimtime="00:02:05.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197440" lastname="AVDIC" firstname="Iman" gender="F" birthdate="2007-09-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.42" eventid="43" heat="2" lane="4">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:04:12.24" eventid="1" heat="2" lane="7">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:04:46.90" eventid="36" heat="2" lane="7">
                  <MEETINFO date="2021-10-31" />
                </ENTRY>
                <ENTRY entrytime="00:08:38.73" eventid="12" heat="2" lane="8">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="25" lane="4" heat="2" heatid="20043" swimtime="00:02:02.30" reactiontime="+67" points="733">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                    <SPLIT distance="75" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:00:58.58" />
                    <SPLIT distance="125" swimtime="00:01:14.31" />
                    <SPLIT distance="150" swimtime="00:01:30.23" />
                    <SPLIT distance="175" swimtime="00:01:46.48" />
                    <SPLIT distance="200" swimtime="00:02:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="24" lane="7" heat="2" heatid="20001" swimtime="00:04:21.65" reactiontime="+71" points="714">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="75" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:00:59.85" />
                    <SPLIT distance="125" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:31.74" />
                    <SPLIT distance="175" swimtime="00:01:47.71" />
                    <SPLIT distance="200" swimtime="00:02:04.29" />
                    <SPLIT distance="225" swimtime="00:02:20.71" />
                    <SPLIT distance="250" swimtime="00:02:37.79" />
                    <SPLIT distance="275" swimtime="00:02:55.03" />
                    <SPLIT distance="300" swimtime="00:03:12.94" />
                    <SPLIT distance="325" swimtime="00:03:30.18" />
                    <SPLIT distance="350" swimtime="00:03:47.65" />
                    <SPLIT distance="375" swimtime="00:04:04.87" />
                    <SPLIT distance="400" swimtime="00:04:21.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="17" lane="7" heat="2" heatid="20036" swimtime="00:04:42.56" reactiontime="+71" points="769">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:47.37" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="125" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:01:42.07" />
                    <SPLIT distance="175" swimtime="00:02:00.14" />
                    <SPLIT distance="200" swimtime="00:02:18.16" />
                    <SPLIT distance="225" swimtime="00:02:38.07" />
                    <SPLIT distance="250" swimtime="00:02:58.10" />
                    <SPLIT distance="275" swimtime="00:03:19.03" />
                    <SPLIT distance="300" swimtime="00:03:39.52" />
                    <SPLIT distance="325" swimtime="00:03:55.99" />
                    <SPLIT distance="350" swimtime="00:04:12.01" />
                    <SPLIT distance="375" swimtime="00:04:27.32" />
                    <SPLIT distance="400" swimtime="00:04:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="18" lane="8" heat="2" heatid="20012" swimtime="00:08:58.28" reactiontime="+71" points="706">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="75" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:01.15" />
                    <SPLIT distance="125" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:33.56" />
                    <SPLIT distance="175" swimtime="00:01:50.33" />
                    <SPLIT distance="200" swimtime="00:02:07.56" />
                    <SPLIT distance="225" swimtime="00:02:24.33" />
                    <SPLIT distance="250" swimtime="00:02:41.28" />
                    <SPLIT distance="275" swimtime="00:02:58.48" />
                    <SPLIT distance="300" swimtime="00:03:15.80" />
                    <SPLIT distance="325" swimtime="00:03:33.07" />
                    <SPLIT distance="350" swimtime="00:03:50.38" />
                    <SPLIT distance="375" swimtime="00:04:07.52" />
                    <SPLIT distance="400" swimtime="00:04:25.06" />
                    <SPLIT distance="425" swimtime="00:04:42.44" />
                    <SPLIT distance="450" swimtime="00:05:00.02" />
                    <SPLIT distance="475" swimtime="00:05:17.09" />
                    <SPLIT distance="500" swimtime="00:05:33.98" />
                    <SPLIT distance="525" swimtime="00:05:51.17" />
                    <SPLIT distance="550" swimtime="00:06:08.72" />
                    <SPLIT distance="575" swimtime="00:06:25.63" />
                    <SPLIT distance="600" swimtime="00:06:42.89" />
                    <SPLIT distance="625" swimtime="00:07:00.28" />
                    <SPLIT distance="650" swimtime="00:07:17.80" />
                    <SPLIT distance="675" swimtime="00:07:34.89" />
                    <SPLIT distance="700" swimtime="00:07:51.95" />
                    <SPLIT distance="725" swimtime="00:08:08.94" />
                    <SPLIT distance="750" swimtime="00:08:25.57" />
                    <SPLIT distance="775" swimtime="00:08:42.18" />
                    <SPLIT distance="800" swimtime="00:08:58.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Belarus" shortname="BLR" code="BLR" nation="BLR" type="NOC">
          <ATHLETES />
        </CLUB>
        <CLUB name="Bolivia" shortname="BOL" code="BOL" nation="BOL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="183473" lastname="NUÑEZ DEL PRADO" firstname="Esteban" gender="M" birthdate="2004-06-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.13" eventid="14" heat="5" lane="2">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.04" eventid="7" heat="2" lane="8">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="57" lane="2" heat="5" heatid="50014" swimtime="00:00:50.76" reactiontime="+61" points="689">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:24.28" />
                    <SPLIT distance="75" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:00:50.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="33" lane="8" heat="2" heatid="20007" swimtime="00:02:01.44" reactiontime="+64" points="735">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                    <SPLIT distance="75" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:00:56.27" />
                    <SPLIT distance="125" swimtime="00:01:13.65" />
                    <SPLIT distance="150" swimtime="00:01:31.66" />
                    <SPLIT distance="175" swimtime="00:01:47.07" />
                    <SPLIT distance="200" swimtime="00:02:01.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124415" lastname="CABRERA" firstname="Jesus" gender="M" birthdate="1997-06-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.50" eventid="41" heat="3" lane="7">
                  <MEETINFO date="2021-08-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="50" lane="7" heat="3" heatid="30041" swimtime="00:00:29.25" reactiontime="+65" points="620">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102175" lastname="TORREZ" firstname="Karen" gender="F" birthdate="1992-07-29">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.66" eventid="13" heat="4" lane="2">
                  <MEETINFO date="2022-10-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.77" eventid="30" heat="5" lane="8">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="42" lane="2" heat="4" heatid="40013" swimtime="00:00:57.19" reactiontime="+61" points="678">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.05" />
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                    <SPLIT distance="75" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:00:57.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="33" lane="8" heat="5" heatid="50030" swimtime="00:00:26.09" reactiontime="+58" points="678">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Botswana" shortname="BOT" code="BOT" nation="BOT" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="145907" lastname="ROBINSON" firstname="Adrian" gender="M" birthdate="2000-04-11">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.57" eventid="16" heat="3" lane="8">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.99" eventid="41" heat="4" lane="3">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="45" lane="8" heat="3" heatid="30016" swimtime="00:01:00.90" reactiontime="+58" points="747">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                    <SPLIT distance="75" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="41" lane="3" heat="4" heatid="40041" swimtime="00:00:27.79" reactiontime="+58" points="723">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.61" />
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129276" lastname="FREEMAN" firstname="James" gender="M" birthdate="2001-03-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.37" eventid="14" heat="5" lane="1">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.63" eventid="44" heat="2" lane="8">
                  <MEETINFO date="2022-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="60" lane="1" heat="5" heatid="50014" swimtime="00:00:51.08" reactiontime="+75" points="676">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.64" />
                    <SPLIT distance="50" swimtime="00:00:24.48" />
                    <SPLIT distance="75" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:00:51.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="39" lane="8" heat="2" heatid="20044" swimtime="00:01:51.02" reactiontime="+71" points="717">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                    <SPLIT distance="75" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:00:54.17" />
                    <SPLIT distance="125" swimtime="00:01:08.14" />
                    <SPLIT distance="150" swimtime="00:01:22.53" />
                    <SPLIT distance="175" swimtime="00:01:37.13" />
                    <SPLIT distance="200" swimtime="00:01:51.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198078" lastname="HUGHES" firstname="Naya" gender="F" birthdate="2004-06-02">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="2" heat="1" lane="6" />
                <ENTRY entrytime="NT" eventid="18" heat="2" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="44" lane="6" heat="1" heatid="10002" swimtime="00:01:09.68" reactiontime="+60" points="488">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="75" swimtime="00:00:51.27" />
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="43" lane="1" heat="2" heatid="20018" swimtime="00:00:32.20" reactiontime="+70" points="483">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Brazil" shortname="BRA" code="BRA" nation="BRA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="124410" lastname="PUMPUTIS" firstname="Caio" gender="M" birthdate="1999-01-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.04" eventid="16" heat="7" lane="6">
                  <MEETINFO date="2021-08-10" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.33" eventid="29" heat="3" lane="5">
                  <MEETINFO date="2021-08-14" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.02" eventid="7" heat="4" lane="6">
                  <MEETINFO date="2021-08-11" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.99" eventid="23" heat="3" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="15" lane="6" heat="7" heatid="70016" swimtime="00:00:57.78" reactiontime="+66" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.66" />
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="75" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:00:57.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="11" lane="8" heat="2" heatid="20216" swimtime="00:00:57.59" reactiontime="+64" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                    <SPLIT distance="75" swimtime="00:00:42.00" />
                    <SPLIT distance="100" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="129" place="-1" lane="8" heat="1" heatid="10129" swimtime="00:02:06.04" status="DSQ" reactiontime="+68" />
                <RESULT eventid="29" place="8" lane="5" heat="3" heatid="30029" swimtime="00:02:04.37" reactiontime="+67" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="75" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:00.48" />
                    <SPLIT distance="125" swimtime="00:01:16.17" />
                    <SPLIT distance="150" swimtime="00:01:32.25" />
                    <SPLIT distance="175" swimtime="00:01:48.00" />
                    <SPLIT distance="200" swimtime="00:02:04.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="15" lane="6" heat="4" heatid="40007" swimtime="00:01:54.65" reactiontime="+66" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:24.42" />
                    <SPLIT distance="75" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:00:53.13" />
                    <SPLIT distance="125" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:26.29" />
                    <SPLIT distance="175" swimtime="00:01:41.13" />
                    <SPLIT distance="200" swimtime="00:01:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="11" lane="3" heat="3" heatid="30023" swimtime="00:00:52.50" reactiontime="+64" points="827">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.05" />
                    <SPLIT distance="50" swimtime="00:00:24.16" />
                    <SPLIT distance="75" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="11" lane="7" heat="2" heatid="20223" swimtime="00:00:52.12" reactiontime="+67" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.64" />
                    <SPLIT distance="50" swimtime="00:00:23.73" />
                    <SPLIT distance="75" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:00:52.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155043" lastname="COELHO SANTOS" firstname="Leonardo" gender="M" birthdate="1995-04-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.53" eventid="39" heat="6" lane="8">
                  <MEETINFO date="2021-08-10" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.50" eventid="7" heat="4" lane="3">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
                <ENTRY entrytime="00:04:06.58" eventid="37" heat="3" lane="2">
                  <MEETINFO date="2021-09-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:52.13" eventid="23" heat="4" lane="6">
                  <MEETINFO date="2021-09-10" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="23" lane="8" heat="6" heatid="60039" swimtime="00:00:51.35" reactiontime="+68" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.94" />
                    <SPLIT distance="50" swimtime="00:00:23.93" />
                    <SPLIT distance="75" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:00:51.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="9" lane="3" heat="4" heatid="40007" swimtime="00:01:53.07" reactiontime="+70" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:24.28" />
                    <SPLIT distance="75" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:00:51.96" />
                    <SPLIT distance="125" swimtime="00:01:08.23" />
                    <SPLIT distance="150" swimtime="00:01:25.29" />
                    <SPLIT distance="175" swimtime="00:01:39.65" />
                    <SPLIT distance="200" swimtime="00:01:53.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="-1" lane="2" heat="3" heatid="30037" swimtime="NT" status="DNS" />
                <RESULT eventid="23" place="12" lane="6" heat="4" heatid="40023" swimtime="00:00:52.58" reactiontime="+69" points="823">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.75" />
                    <SPLIT distance="50" swimtime="00:00:23.61" />
                    <SPLIT distance="75" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:00:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="13" lane="7" heat="1" heatid="10223" swimtime="00:00:52.37" reactiontime="+68" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.80" />
                    <SPLIT distance="50" swimtime="00:00:23.56" />
                    <SPLIT distance="75" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124426" lastname="SPAJARI" firstname="Pedro" gender="M" birthdate="1997-02-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.70" eventid="14" heat="11" lane="6">
                  <MEETINFO date="2021-09-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.41" eventid="31" heat="8" lane="4">
                  <MEETINFO date="2021-09-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="14" lane="6" heat="11" heatid="110014" swimtime="00:00:46.94" reactiontime="+62" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.79" />
                    <SPLIT distance="50" swimtime="00:00:22.67" />
                    <SPLIT distance="75" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:00:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="16" lane="1" heat="1" heatid="10214" swimtime="00:00:47.32" reactiontime="+64" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.48" />
                    <SPLIT distance="75" swimtime="00:00:34.85" />
                    <SPLIT distance="100" swimtime="00:00:47.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="42" lane="4" heat="8" heatid="80031" swimtime="00:00:21.84" reactiontime="+62" points="786">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.59" />
                    <SPLIT distance="50" swimtime="00:00:21.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144007" lastname="SANTOS" firstname="Gabriel" gender="M" birthdate="1996-05-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.39" eventid="14" heat="10" lane="3">
                  <MEETINFO date="2022-09-15" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.40" eventid="5" heat="6" lane="3">
                  <MEETINFO date="2022-04-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="23" lane="3" heat="10" heatid="100014" swimtime="00:00:47.14" reactiontime="+59" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.66" />
                    <SPLIT distance="50" swimtime="00:00:22.65" />
                    <SPLIT distance="75" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:00:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="25" lane="3" heat="6" heatid="60005" swimtime="00:00:22.89" reactiontime="+58" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.28" />
                    <SPLIT distance="50" swimtime="00:00:22.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143708" lastname="CORREIA" firstname="Breno" gender="M" birthdate="1999-02-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.80" eventid="44" heat="4" lane="2">
                  <MEETINFO date="2022-09-16" />
                </ENTRY>
                <ENTRY entrytime="00:03:42.42" eventid="24" heat="3" lane="4">
                  <MEETINFO date="2022-08-10" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="14" lane="2" heat="4" heatid="40044" swimtime="00:01:43.48" reactiontime="+58" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:24.26" />
                    <SPLIT distance="75" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:00:50.68" />
                    <SPLIT distance="125" swimtime="00:01:03.89" />
                    <SPLIT distance="150" swimtime="00:01:17.13" />
                    <SPLIT distance="175" swimtime="00:01:30.50" />
                    <SPLIT distance="200" swimtime="00:01:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="13" lane="4" heat="3" heatid="30024" swimtime="00:03:41.89" reactiontime="+61" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                    <SPLIT distance="75" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:00:53.24" />
                    <SPLIT distance="125" swimtime="00:01:07.33" />
                    <SPLIT distance="150" swimtime="00:01:21.28" />
                    <SPLIT distance="175" swimtime="00:01:35.56" />
                    <SPLIT distance="200" swimtime="00:01:49.67" />
                    <SPLIT distance="225" swimtime="00:02:03.97" />
                    <SPLIT distance="250" swimtime="00:02:18.18" />
                    <SPLIT distance="275" swimtime="00:02:32.57" />
                    <SPLIT distance="300" swimtime="00:02:46.78" />
                    <SPLIT distance="325" swimtime="00:03:00.97" />
                    <SPLIT distance="350" swimtime="00:03:15.00" />
                    <SPLIT distance="375" swimtime="00:03:28.77" />
                    <SPLIT distance="400" swimtime="00:03:41.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101084" lastname="GOMES JUNIOR" firstname="Joao" gender="M" birthdate="1986-01-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.80" eventid="41" heat="8" lane="5">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="-1" lane="5" heat="8" heatid="80041" swimtime="00:00:26.20" status="DSQ" reactiontime="+67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101178" lastname="SANTOS" firstname="Nicholas" gender="M" birthdate="1980-02-14">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.81" eventid="5" heat="9" lane="4">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="105" place="1" lane="6" heat="1" heatid="10105" swimtime="00:00:21.78" reactiontime="+60" points="995">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.00" />
                    <SPLIT distance="50" swimtime="00:00:21.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="14" lane="4" heat="9" heatid="90005" swimtime="00:00:22.46" reactiontime="+60" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.15" />
                    <SPLIT distance="50" swimtime="00:00:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="4" lane="1" heat="1" heatid="10205" swimtime="00:00:22.08" reactiontime="+61" points="955">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.02" />
                    <SPLIT distance="50" swimtime="00:00:22.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110357" lastname="TOMANIK DIAMANTE" firstname="Giovanna" gender="F" birthdate="1997-06-26">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:56.79" eventid="38" heat="4" lane="6">
                  <MEETINFO date="2022-08-10" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.15" eventid="20" heat="3" lane="2">
                  <MEETINFO date="2022-09-15" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.05" eventid="43" heat="3" lane="6">
                  <MEETINFO date="2022-09-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:00:26.19" eventid="4" heat="4" lane="7">
                  <MEETINFO date="2022-09-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="14" lane="6" heat="4" heatid="40038" swimtime="00:00:57.50" reactiontime="+66" points="855">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                    <SPLIT distance="75" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:00:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="12" lane="1" heat="1" heatid="10238" swimtime="00:00:57.13" reactiontime="+64" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                    <SPLIT distance="75" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:00:57.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="16" lane="2" heat="3" heatid="30020" swimtime="00:02:09.60" reactiontime="+67" points="786">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.36" />
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                    <SPLIT distance="75" swimtime="00:00:45.27" />
                    <SPLIT distance="100" swimtime="00:01:01.37" />
                    <SPLIT distance="125" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:01:34.23" />
                    <SPLIT distance="175" swimtime="00:01:51.66" />
                    <SPLIT distance="200" swimtime="00:02:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="18" lane="6" heat="3" heatid="30043" swimtime="00:01:57.44" reactiontime="+64" points="828">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.02" />
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                    <SPLIT distance="75" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:00:56.72" />
                    <SPLIT distance="125" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:26.63" />
                    <SPLIT distance="175" swimtime="00:01:42.04" />
                    <SPLIT distance="200" swimtime="00:01:57.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="26" lane="7" heat="4" heatid="40004" swimtime="00:00:26.48" reactiontime="+67" points="780">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202143" lastname="BALDUCCINI" firstname="Stephanie" gender="F" birthdate="2004-09-20">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:53.36" eventid="13" heat="9" lane="1">
                  <MEETINFO date="2022-09-15" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.02" eventid="43" heat="4" lane="6">
                  <MEETINFO date="2022-09-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.99" eventid="6" heat="5" lane="8">
                  <MEETINFO date="2021-08-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:00:24.97" eventid="30" heat="7" lane="8">
                  <MEETINFO date="2021-08-14" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.84" eventid="22" heat="4" lane="1">
                  <MEETINFO date="2021-08-14" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="16" lane="1" heat="9" heatid="90013" swimtime="00:00:53.32" reactiontime="+65" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.44" />
                    <SPLIT distance="50" swimtime="00:00:25.94" />
                    <SPLIT distance="75" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:00:53.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="16" lane="8" heat="1" heatid="10213" swimtime="00:00:53.64" reactiontime="+72" points="822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:25.92" />
                    <SPLIT distance="75" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="16" lane="6" heat="4" heatid="40043" swimtime="00:01:57.09" reactiontime="+69" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="75" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:00:57.23" />
                    <SPLIT distance="125" swimtime="00:01:12.12" />
                    <SPLIT distance="150" swimtime="00:01:27.05" />
                    <SPLIT distance="175" swimtime="00:01:42.42" />
                    <SPLIT distance="200" swimtime="00:01:57.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="25" lane="8" heat="5" heatid="50006" swimtime="00:02:12.46" reactiontime="+69" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:45.06" />
                    <SPLIT distance="100" swimtime="00:01:01.10" />
                    <SPLIT distance="125" swimtime="00:01:20.42" />
                    <SPLIT distance="150" swimtime="00:01:40.62" />
                    <SPLIT distance="175" swimtime="00:01:57.21" />
                    <SPLIT distance="200" swimtime="00:02:12.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="28" lane="8" heat="7" heatid="70030" swimtime="00:00:25.24" reactiontime="+70" points="749">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="20" lane="1" heat="4" heatid="40022" swimtime="00:01:01.58" reactiontime="+71" points="772">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="75" swimtime="00:00:46.69" />
                    <SPLIT distance="100" swimtime="00:01:01.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108174" lastname="RONCATTO" firstname="Gabrielle" gender="F" birthdate="1998-07-19">
              <ENTRIES>
                <ENTRY entrytime="00:04:03.77" eventid="1" heat="4" lane="1">
                  <MEETINFO date="2022-08-10" />
                </ENTRY>
                <ENTRY entrytime="00:04:36.38" eventid="36" heat="4" lane="8">
                  <MEETINFO date="2022-09-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:08:26.37" eventid="12" heat="2" lane="3">
                  <MEETINFO date="2022-09-14" />
                </ENTRY>
                <ENTRY entrytime="00:15:56.09" eventid="33" heat="0" lane="2147483647">
                  <MEETINFO date="2022-09-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="13" lane="1" heat="4" heatid="40001" swimtime="00:04:08.39" reactiontime="+71" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:00:57.67" />
                    <SPLIT distance="125" swimtime="00:01:12.88" />
                    <SPLIT distance="150" swimtime="00:01:28.35" />
                    <SPLIT distance="175" swimtime="00:01:43.86" />
                    <SPLIT distance="200" swimtime="00:01:59.80" />
                    <SPLIT distance="225" swimtime="00:02:15.70" />
                    <SPLIT distance="250" swimtime="00:02:31.67" />
                    <SPLIT distance="275" swimtime="00:02:47.81" />
                    <SPLIT distance="300" swimtime="00:03:03.95" />
                    <SPLIT distance="325" swimtime="00:03:20.26" />
                    <SPLIT distance="350" swimtime="00:03:36.62" />
                    <SPLIT distance="375" swimtime="00:03:53.00" />
                    <SPLIT distance="400" swimtime="00:04:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="-1" lane="8" heat="4" heatid="40036" swimtime="NT" status="DNS" />
                <RESULT eventid="112" place="8" lane="3" heat="2" heatid="20012" swimtime="00:08:25.45" reactiontime="+73" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="75" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:00.40" />
                    <SPLIT distance="125" swimtime="00:01:16.30" />
                    <SPLIT distance="150" swimtime="00:01:32.16" />
                    <SPLIT distance="175" swimtime="00:01:48.02" />
                    <SPLIT distance="200" swimtime="00:02:04.08" />
                    <SPLIT distance="225" swimtime="00:02:20.08" />
                    <SPLIT distance="250" swimtime="00:02:35.99" />
                    <SPLIT distance="275" swimtime="00:02:51.95" />
                    <SPLIT distance="300" swimtime="00:03:07.98" />
                    <SPLIT distance="325" swimtime="00:03:24.02" />
                    <SPLIT distance="350" swimtime="00:03:40.03" />
                    <SPLIT distance="375" swimtime="00:03:55.95" />
                    <SPLIT distance="400" swimtime="00:04:12.05" />
                    <SPLIT distance="425" swimtime="00:04:27.98" />
                    <SPLIT distance="450" swimtime="00:04:43.95" />
                    <SPLIT distance="475" swimtime="00:04:59.92" />
                    <SPLIT distance="500" swimtime="00:05:15.81" />
                    <SPLIT distance="525" swimtime="00:05:31.75" />
                    <SPLIT distance="550" swimtime="00:05:47.71" />
                    <SPLIT distance="575" swimtime="00:06:03.65" />
                    <SPLIT distance="600" swimtime="00:06:19.56" />
                    <SPLIT distance="625" swimtime="00:06:35.56" />
                    <SPLIT distance="650" swimtime="00:06:51.54" />
                    <SPLIT distance="675" swimtime="00:07:07.56" />
                    <SPLIT distance="700" swimtime="00:07:23.54" />
                    <SPLIT distance="725" swimtime="00:07:39.52" />
                    <SPLIT distance="750" swimtime="00:07:55.38" />
                    <SPLIT distance="775" swimtime="00:08:11.21" />
                    <SPLIT distance="800" swimtime="00:08:25.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="12" lane="2" heat="5" heatid="30133" swimtime="00:16:33.31" reactiontime="+70" points="789">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                    <SPLIT distance="75" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="125" swimtime="00:01:15.71" />
                    <SPLIT distance="150" swimtime="00:01:31.67" />
                    <SPLIT distance="175" swimtime="00:01:47.73" />
                    <SPLIT distance="200" swimtime="00:02:03.56" />
                    <SPLIT distance="225" swimtime="00:02:19.49" />
                    <SPLIT distance="250" swimtime="00:02:35.49" />
                    <SPLIT distance="275" swimtime="00:02:51.57" />
                    <SPLIT distance="300" swimtime="00:03:07.59" />
                    <SPLIT distance="325" swimtime="00:03:23.61" />
                    <SPLIT distance="350" swimtime="00:03:39.69" />
                    <SPLIT distance="375" swimtime="00:03:55.62" />
                    <SPLIT distance="400" swimtime="00:04:11.67" />
                    <SPLIT distance="425" swimtime="00:04:27.69" />
                    <SPLIT distance="450" swimtime="00:04:43.80" />
                    <SPLIT distance="475" swimtime="00:04:59.93" />
                    <SPLIT distance="500" swimtime="00:05:16.11" />
                    <SPLIT distance="525" swimtime="00:05:32.26" />
                    <SPLIT distance="550" swimtime="00:05:48.78" />
                    <SPLIT distance="575" swimtime="00:06:05.09" />
                    <SPLIT distance="600" swimtime="00:06:21.42" />
                    <SPLIT distance="625" swimtime="00:06:37.79" />
                    <SPLIT distance="650" swimtime="00:06:54.52" />
                    <SPLIT distance="675" swimtime="00:07:10.99" />
                    <SPLIT distance="700" swimtime="00:07:27.52" />
                    <SPLIT distance="725" swimtime="00:07:44.24" />
                    <SPLIT distance="750" swimtime="00:08:00.76" />
                    <SPLIT distance="775" swimtime="00:08:17.55" />
                    <SPLIT distance="800" swimtime="00:08:34.24" />
                    <SPLIT distance="825" swimtime="00:08:50.83" />
                    <SPLIT distance="850" swimtime="00:09:07.67" />
                    <SPLIT distance="875" swimtime="00:09:24.57" />
                    <SPLIT distance="900" swimtime="00:09:41.60" />
                    <SPLIT distance="925" swimtime="00:09:58.60" />
                    <SPLIT distance="950" swimtime="00:10:15.59" />
                    <SPLIT distance="975" swimtime="00:10:32.72" />
                    <SPLIT distance="1000" swimtime="00:10:49.95" />
                    <SPLIT distance="1025" swimtime="00:11:07.07" />
                    <SPLIT distance="1050" swimtime="00:11:24.43" />
                    <SPLIT distance="1075" swimtime="00:11:41.69" />
                    <SPLIT distance="1100" swimtime="00:11:59.04" />
                    <SPLIT distance="1125" swimtime="00:12:16.25" />
                    <SPLIT distance="1150" swimtime="00:12:33.79" />
                    <SPLIT distance="1175" swimtime="00:12:51.10" />
                    <SPLIT distance="1200" swimtime="00:13:08.67" />
                    <SPLIT distance="1225" swimtime="00:13:25.97" />
                    <SPLIT distance="1250" swimtime="00:13:43.39" />
                    <SPLIT distance="1275" swimtime="00:14:00.49" />
                    <SPLIT distance="1300" swimtime="00:14:17.58" />
                    <SPLIT distance="1325" swimtime="00:14:34.80" />
                    <SPLIT distance="1350" swimtime="00:14:52.01" />
                    <SPLIT distance="1375" swimtime="00:15:09.03" />
                    <SPLIT distance="1400" swimtime="00:15:26.17" />
                    <SPLIT distance="1425" swimtime="00:15:43.15" />
                    <SPLIT distance="1450" swimtime="00:16:00.30" />
                    <SPLIT distance="1475" swimtime="00:16:17.11" />
                    <SPLIT distance="1500" swimtime="00:16:33.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143700" lastname="PEIXOTO" firstname="Lucas" gender="M" birthdate="2000-09-05" />
            <ATHLETE athleteid="202142" lastname="RODRIGUES" firstname="Aline" gender="F" birthdate="1995-04-07" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Brazil">
              <RESULTS>
                <RESULT eventid="109" place="4" lane="5" heat="1" swimtime="00:03:06.85" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:22.23" />
                    <SPLIT distance="75" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:00:47.04" />
                    <SPLIT distance="125" swimtime="00:00:57.51" />
                    <SPLIT distance="150" swimtime="00:01:09.33" />
                    <SPLIT distance="175" swimtime="00:01:21.58" />
                    <SPLIT distance="200" swimtime="00:01:33.68" />
                    <SPLIT distance="225" swimtime="00:01:43.95" />
                    <SPLIT distance="250" swimtime="00:01:55.64" />
                    <SPLIT distance="275" swimtime="00:02:07.91" />
                    <SPLIT distance="300" swimtime="00:02:20.22" />
                    <SPLIT distance="325" swimtime="00:02:30.56" />
                    <SPLIT distance="350" swimtime="00:02:42.21" />
                    <SPLIT distance="375" swimtime="00:02:54.70" />
                    <SPLIT distance="400" swimtime="00:03:06.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="144007" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="143708" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="143700" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="124426" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="2" lane="5" heat="1" swimtime="00:03:06.82" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.47" />
                    <SPLIT distance="50" swimtime="00:00:22.52" />
                    <SPLIT distance="75" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:00:47.31" />
                    <SPLIT distance="125" swimtime="00:00:57.73" />
                    <SPLIT distance="150" swimtime="00:01:09.38" />
                    <SPLIT distance="175" swimtime="00:01:21.33" />
                    <SPLIT distance="200" swimtime="00:01:33.27" />
                    <SPLIT distance="225" swimtime="00:01:43.31" />
                    <SPLIT distance="250" swimtime="00:01:55.24" />
                    <SPLIT distance="275" swimtime="00:02:07.50" />
                    <SPLIT distance="300" swimtime="00:02:20.03" />
                    <SPLIT distance="325" swimtime="00:02:30.38" />
                    <SPLIT distance="350" swimtime="00:02:42.37" />
                    <SPLIT distance="375" swimtime="00:02:54.54" />
                    <SPLIT distance="400" swimtime="00:03:06.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="144007" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="143708" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="143700" reactiontime="+6" />
                    <RELAYPOSITION number="4" athleteid="124426" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Brazil">
              <RESULTS>
                <RESULT eventid="48" place="-1" lane="5" heat="3" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Brazil">
              <RESULTS>
                <RESULT eventid="32" place="9" lane="4" heat="1" swimtime="00:07:02.32" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:24.25" />
                    <SPLIT distance="75" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:00:50.85" />
                    <SPLIT distance="125" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:17.91" />
                    <SPLIT distance="175" swimtime="00:01:31.75" />
                    <SPLIT distance="200" swimtime="00:01:45.45" />
                    <SPLIT distance="225" swimtime="00:01:56.47" />
                    <SPLIT distance="250" swimtime="00:02:09.16" />
                    <SPLIT distance="275" swimtime="00:02:22.27" />
                    <SPLIT distance="300" swimtime="00:02:35.67" />
                    <SPLIT distance="325" swimtime="00:02:49.21" />
                    <SPLIT distance="350" swimtime="00:03:02.77" />
                    <SPLIT distance="375" swimtime="00:03:16.17" />
                    <SPLIT distance="400" swimtime="00:03:28.97" />
                    <SPLIT distance="425" swimtime="00:03:39.69" />
                    <SPLIT distance="450" swimtime="00:03:52.49" />
                    <SPLIT distance="475" swimtime="00:04:05.79" />
                    <SPLIT distance="500" swimtime="00:04:19.23" />
                    <SPLIT distance="525" swimtime="00:04:32.92" />
                    <SPLIT distance="550" swimtime="00:04:46.70" />
                    <SPLIT distance="575" swimtime="00:05:00.48" />
                    <SPLIT distance="600" swimtime="00:05:13.85" />
                    <SPLIT distance="625" swimtime="00:05:24.95" />
                    <SPLIT distance="650" swimtime="00:05:37.77" />
                    <SPLIT distance="675" swimtime="00:05:50.97" />
                    <SPLIT distance="700" swimtime="00:06:04.62" />
                    <SPLIT distance="725" swimtime="00:06:18.61" />
                    <SPLIT distance="750" swimtime="00:06:33.03" />
                    <SPLIT distance="775" swimtime="00:06:47.75" />
                    <SPLIT distance="800" swimtime="00:07:02.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="143700" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="143708" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="155043" reactiontime="+22" />
                    <RELAYPOSITION number="4" athleteid="124426" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Brazil">
              <RESULTS>
                <RESULT eventid="126" place="8" lane="7" heat="1" swimtime="00:01:26.34" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.42" />
                    <SPLIT distance="50" swimtime="00:00:21.77" />
                    <SPLIT distance="75" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:00:43.58" />
                    <SPLIT distance="125" swimtime="00:00:53.48" />
                    <SPLIT distance="150" swimtime="00:01:05.21" />
                    <SPLIT distance="175" swimtime="00:01:15.16" />
                    <SPLIT distance="200" swimtime="00:01:26.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124426" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="144007" reactiontime="+27" />
                    <RELAYPOSITION number="3" athleteid="101178" reactiontime="+12" />
                    <RELAYPOSITION number="4" athleteid="143700" reactiontime="+12" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="6" lane="6" heat="2" swimtime="00:01:26.10" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.38" />
                    <SPLIT distance="50" swimtime="00:00:21.79" />
                    <SPLIT distance="75" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:00:43.10" />
                    <SPLIT distance="125" swimtime="00:00:53.09" />
                    <SPLIT distance="150" swimtime="00:01:04.77" />
                    <SPLIT distance="175" swimtime="00:01:14.79" />
                    <SPLIT distance="200" swimtime="00:01:26.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="144007" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="124426" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="101178" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="143700" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Brazil">
              <RESULTS>
                <RESULT eventid="127" place="8" lane="8" heat="1" swimtime="00:01:32.17" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.57" />
                    <SPLIT distance="50" swimtime="00:00:21.85" />
                    <SPLIT distance="75" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:00:43.02" />
                    <SPLIT distance="125" swimtime="00:00:55.04" />
                    <SPLIT distance="150" swimtime="00:01:07.85" />
                    <SPLIT distance="175" swimtime="00:01:19.52" />
                    <SPLIT distance="200" swimtime="00:01:32.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="143700" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="124426" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="202143" reactiontime="+16" />
                    <RELAYPOSITION number="4" athleteid="110357" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="8" lane="8" heat="2" swimtime="00:01:32.15" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.49" />
                    <SPLIT distance="50" swimtime="00:00:21.73" />
                    <SPLIT distance="75" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:00:43.13" />
                    <SPLIT distance="125" swimtime="00:00:54.79" />
                    <SPLIT distance="150" swimtime="00:01:07.46" />
                    <SPLIT distance="175" swimtime="00:01:19.44" />
                    <SPLIT distance="200" swimtime="00:01:32.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="143700" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="124426" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="202143" reactiontime="+6" />
                    <RELAYPOSITION number="4" athleteid="110357" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Brazil">
              <RESULTS>
                <RESULT eventid="8" place="9" lane="2" heat="2" swimtime="00:03:38.61" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                    <SPLIT distance="75" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:00:53.99" />
                    <SPLIT distance="125" swimtime="00:01:06.54" />
                    <SPLIT distance="150" swimtime="00:01:20.29" />
                    <SPLIT distance="175" swimtime="00:01:34.17" />
                    <SPLIT distance="200" swimtime="00:01:47.81" />
                    <SPLIT distance="225" swimtime="00:02:00.30" />
                    <SPLIT distance="250" swimtime="00:02:14.21" />
                    <SPLIT distance="275" swimtime="00:02:28.57" />
                    <SPLIT distance="300" swimtime="00:02:42.89" />
                    <SPLIT distance="325" swimtime="00:02:55.94" />
                    <SPLIT distance="350" swimtime="00:03:10.06" />
                    <SPLIT distance="375" swimtime="00:03:24.63" />
                    <SPLIT distance="400" swimtime="00:03:38.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="110357" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="202143" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="202142" reactiontime="+47" />
                    <RELAYPOSITION number="4" athleteid="108174" reactiontime="+55" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Brazil">
              <RESULTS>
                <RESULT eventid="117" place="7" lane="7" heat="1" swimtime="00:07:48.83" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                    <SPLIT distance="75" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:00:57.20" />
                    <SPLIT distance="125" swimtime="00:01:12.14" />
                    <SPLIT distance="150" swimtime="00:01:27.46" />
                    <SPLIT distance="175" swimtime="00:01:42.91" />
                    <SPLIT distance="200" swimtime="00:01:58.05" />
                    <SPLIT distance="225" swimtime="00:02:10.62" />
                    <SPLIT distance="250" swimtime="00:02:24.80" />
                    <SPLIT distance="275" swimtime="00:02:39.11" />
                    <SPLIT distance="300" swimtime="00:02:53.61" />
                    <SPLIT distance="325" swimtime="00:03:08.33" />
                    <SPLIT distance="350" swimtime="00:03:23.58" />
                    <SPLIT distance="375" swimtime="00:03:39.26" />
                    <SPLIT distance="400" swimtime="00:03:54.64" />
                    <SPLIT distance="425" swimtime="00:04:07.38" />
                    <SPLIT distance="450" swimtime="00:04:21.48" />
                    <SPLIT distance="475" swimtime="00:04:36.01" />
                    <SPLIT distance="500" swimtime="00:04:50.80" />
                    <SPLIT distance="525" swimtime="00:05:05.83" />
                    <SPLIT distance="550" swimtime="00:05:21.12" />
                    <SPLIT distance="575" swimtime="00:05:36.43" />
                    <SPLIT distance="600" swimtime="00:05:51.10" />
                    <SPLIT distance="625" swimtime="00:06:03.92" />
                    <SPLIT distance="650" swimtime="00:06:18.52" />
                    <SPLIT distance="675" swimtime="00:06:33.38" />
                    <SPLIT distance="700" swimtime="00:06:48.42" />
                    <SPLIT distance="725" swimtime="00:07:03.64" />
                    <SPLIT distance="750" swimtime="00:07:18.88" />
                    <SPLIT distance="775" swimtime="00:07:34.27" />
                    <SPLIT distance="800" swimtime="00:07:48.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202143" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="110357" reactiontime="+40" />
                    <RELAYPOSITION number="3" athleteid="108174" reactiontime="+47" />
                    <RELAYPOSITION number="4" athleteid="202142" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="6" lane="3" heat="2" swimtime="00:07:48.42" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.21" />
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="75" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:00:57.23" />
                    <SPLIT distance="125" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:27.04" />
                    <SPLIT distance="175" swimtime="00:01:41.97" />
                    <SPLIT distance="200" swimtime="00:01:56.55" />
                    <SPLIT distance="225" swimtime="00:02:09.15" />
                    <SPLIT distance="250" swimtime="00:02:23.44" />
                    <SPLIT distance="275" swimtime="00:02:38.05" />
                    <SPLIT distance="300" swimtime="00:02:52.85" />
                    <SPLIT distance="325" swimtime="00:03:07.50" />
                    <SPLIT distance="350" swimtime="00:03:22.67" />
                    <SPLIT distance="375" swimtime="00:03:38.07" />
                    <SPLIT distance="400" swimtime="00:03:53.34" />
                    <SPLIT distance="425" swimtime="00:04:06.21" />
                    <SPLIT distance="450" swimtime="00:04:20.65" />
                    <SPLIT distance="475" swimtime="00:04:35.34" />
                    <SPLIT distance="500" swimtime="00:04:50.21" />
                    <SPLIT distance="525" swimtime="00:05:05.29" />
                    <SPLIT distance="550" swimtime="00:05:20.48" />
                    <SPLIT distance="575" swimtime="00:05:35.52" />
                    <SPLIT distance="600" swimtime="00:05:49.91" />
                    <SPLIT distance="625" swimtime="00:06:02.30" />
                    <SPLIT distance="650" swimtime="00:06:16.83" />
                    <SPLIT distance="675" swimtime="00:06:31.43" />
                    <SPLIT distance="700" swimtime="00:06:46.36" />
                    <SPLIT distance="725" swimtime="00:07:01.83" />
                    <SPLIT distance="750" swimtime="00:07:17.33" />
                    <SPLIT distance="775" swimtime="00:07:33.01" />
                    <SPLIT distance="800" swimtime="00:07:48.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202143" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="110357" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="108174" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="202142" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Brazil">
              <RESULTS>
                <RESULT eventid="35" place="-1" lane="6" heat="1" status="DSQ" swimtime="00:01:35.57" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:24.35" />
                    <SPLIT distance="75" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:00:51.04" />
                    <SPLIT distance="125" swimtime="00:01:01.36" />
                    <SPLIT distance="150" swimtime="00:01:14.34" />
                    <SPLIT distance="175" swimtime="00:01:24.48" />
                    <SPLIT distance="200" swimtime="00:01:35.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="155043" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="124410" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="144007" reactiontime="+26" status="DSQ" />
                    <RELAYPOSITION number="4" athleteid="143700" reactiontime="+22" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Bahrain" shortname="BRN" code="BRN" nation="BRN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="213240" lastname="ALOBAIDLI" firstname="Amani" gender="F" birthdate="2006-01-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.74" eventid="2" heat="2" lane="2">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.38" eventid="18" heat="3" lane="4">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="38" lane="2" heat="2" heatid="20002" swimtime="00:01:03.37" reactiontime="+70" points="649">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="75" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:03.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="34" lane="4" heat="3" heatid="30018" swimtime="00:00:28.76" reactiontime="+66" points="678">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.27" />
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Brunei Darussalam" shortname="BRU" code="BRU" nation="BRU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="100454" lastname="AHMAD" firstname="Muhammad Isa" gender="M" birthdate="1998-02-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.09" eventid="16" heat="2" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.32" eventid="41" heat="3" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="55" lane="7" heat="2" heatid="20016" swimtime="00:01:05.15" reactiontime="+68" points="610">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="75" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="-1" lane="2" heat="3" heatid="30041" swimtime="00:00:29.42" status="DSQ" reactiontime="+67" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Bulgaria" shortname="BUL" code="BUL" nation="BUL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="163143" lastname="LEVTEROV" firstname="Kaloyan" gender="M" birthdate="2003-02-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.21" eventid="3" heat="3" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.26" eventid="46" heat="4" lane="8">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="31" lane="6" heat="3" heatid="30003" swimtime="00:00:53.22" reactiontime="+52" points="748">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.61" />
                    <SPLIT distance="50" swimtime="00:00:25.77" />
                    <SPLIT distance="75" swimtime="00:00:39.46" />
                    <SPLIT distance="100" swimtime="00:00:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="21" lane="8" heat="4" heatid="40046" swimtime="00:01:55.98" reactiontime="+54" points="755">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:00:56.54" />
                    <SPLIT distance="125" swimtime="00:01:11.14" />
                    <SPLIT distance="150" swimtime="00:01:25.94" />
                    <SPLIT distance="175" swimtime="00:01:40.91" />
                    <SPLIT distance="200" swimtime="00:01:55.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213077" lastname="SABEV" firstname="Tonislav" gender="M" birthdate="2002-12-13">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.39" eventid="16" heat="3" lane="1">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:27.58" eventid="41" heat="5" lane="1">
                  <MEETINFO date="2022-08-15" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="29" lane="1" heat="3" heatid="30016" swimtime="00:00:58.58" reactiontime="+64" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                    <SPLIT distance="75" swimtime="00:00:42.48" />
                    <SPLIT distance="100" swimtime="00:00:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="-1" lane="1" heat="5" heatid="50041" swimtime="00:00:26.55" status="DSQ" reactiontime="+65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105113" lastname="IVANOV" firstname="Antani" gender="M" birthdate="1999-07-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.20" eventid="39" heat="7" lane="7">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.49" eventid="21" heat="3" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="27" lane="7" heat="7" heatid="70039" swimtime="00:00:51.70" reactiontime="+69" points="789">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.16" />
                    <SPLIT distance="50" swimtime="00:00:24.23" />
                    <SPLIT distance="75" swimtime="00:00:37.77" />
                    <SPLIT distance="100" swimtime="00:00:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="13" lane="6" heat="3" heatid="30021" swimtime="00:01:52.38" reactiontime="+69" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:25.17" />
                    <SPLIT distance="75" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:00:53.38" />
                    <SPLIT distance="125" swimtime="00:01:07.89" />
                    <SPLIT distance="150" swimtime="00:01:22.57" />
                    <SPLIT distance="175" swimtime="00:01:37.61" />
                    <SPLIT distance="200" swimtime="00:01:52.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202468" lastname="NANKOV" firstname="Deniel Genadiev" gender="M" birthdate="2003-01-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.33" eventid="14" heat="6" lane="7">
                  <MEETINFO date="2022-04-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.58" eventid="31" heat="6" lane="1">
                  <MEETINFO date="2022-08-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="25" lane="7" heat="6" heatid="60014" swimtime="00:00:47.30" reactiontime="+62" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.75" />
                    <SPLIT distance="50" swimtime="00:00:22.41" />
                    <SPLIT distance="75" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="44" lane="1" heat="6" heatid="60031" swimtime="00:00:21.89" reactiontime="+61" points="781">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.61" />
                    <SPLIT distance="50" swimtime="00:00:21.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213076" lastname="MITSIN" firstname="Petar Petrov" gender="M" birthdate="2005-08-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:44.36" eventid="44" heat="4" lane="1">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="14" lane="1" heat="4" heatid="40044" swimtime="00:01:43.48" reactiontime="+63" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                    <SPLIT distance="75" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:00:49.99" />
                    <SPLIT distance="125" swimtime="00:01:03.19" />
                    <SPLIT distance="150" swimtime="00:01:16.56" />
                    <SPLIT distance="175" swimtime="00:01:30.29" />
                    <SPLIT distance="200" swimtime="00:01:43.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="142443" lastname="BRATANOV" firstname="Kaloyan" gender="M" birthdate="2000-07-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.28" eventid="7" heat="4" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="14" lane="7" heat="4" heatid="40007" swimtime="00:01:54.50" reactiontime="+69" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.22" />
                    <SPLIT distance="50" swimtime="00:00:24.83" />
                    <SPLIT distance="75" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:00:54.12" />
                    <SPLIT distance="125" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:26.97" />
                    <SPLIT distance="175" swimtime="00:01:41.32" />
                    <SPLIT distance="200" swimtime="00:01:54.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149077" lastname="YANCHEV" firstname="Yordan" gender="M" birthdate="2001-08-30">
              <ENTRIES>
                <ENTRY entrytime="00:03:48.12" eventid="24" heat="2" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:08:15.39" eventid="42" heat="1" lane="7">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="24" place="19" lane="6" heat="2" heatid="20024" swimtime="00:03:45.70" reactiontime="+69" points="831">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                    <SPLIT distance="75" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:00:53.81" />
                    <SPLIT distance="125" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:22.04" />
                    <SPLIT distance="175" swimtime="00:01:36.13" />
                    <SPLIT distance="200" swimtime="00:01:50.54" />
                    <SPLIT distance="225" swimtime="00:02:04.53" />
                    <SPLIT distance="250" swimtime="00:02:18.77" />
                    <SPLIT distance="275" swimtime="00:02:32.90" />
                    <SPLIT distance="300" swimtime="00:02:47.29" />
                    <SPLIT distance="325" swimtime="00:03:01.64" />
                    <SPLIT distance="350" swimtime="00:03:16.34" />
                    <SPLIT distance="375" swimtime="00:03:31.23" />
                    <SPLIT distance="400" swimtime="00:03:45.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="21" lane="7" heat="1" heatid="10042" swimtime="00:08:17.85" reactiontime="+70" points="706">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="75" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:00:57.63" />
                    <SPLIT distance="125" swimtime="00:01:12.59" />
                    <SPLIT distance="150" swimtime="00:01:27.77" />
                    <SPLIT distance="175" swimtime="00:01:42.91" />
                    <SPLIT distance="200" swimtime="00:01:58.20" />
                    <SPLIT distance="225" swimtime="00:02:13.42" />
                    <SPLIT distance="250" swimtime="00:02:28.79" />
                    <SPLIT distance="275" swimtime="00:02:44.14" />
                    <SPLIT distance="300" swimtime="00:02:59.62" />
                    <SPLIT distance="325" swimtime="00:03:15.14" />
                    <SPLIT distance="350" swimtime="00:03:30.64" />
                    <SPLIT distance="375" swimtime="00:03:46.28" />
                    <SPLIT distance="400" swimtime="00:04:02.01" />
                    <SPLIT distance="425" swimtime="00:04:17.46" />
                    <SPLIT distance="450" swimtime="00:04:33.28" />
                    <SPLIT distance="475" swimtime="00:04:49.06" />
                    <SPLIT distance="500" swimtime="00:05:05.06" />
                    <SPLIT distance="525" swimtime="00:05:21.25" />
                    <SPLIT distance="550" swimtime="00:05:37.36" />
                    <SPLIT distance="575" swimtime="00:05:53.56" />
                    <SPLIT distance="600" swimtime="00:06:09.76" />
                    <SPLIT distance="625" swimtime="00:06:25.88" />
                    <SPLIT distance="650" swimtime="00:06:41.87" />
                    <SPLIT distance="675" swimtime="00:06:57.96" />
                    <SPLIT distance="700" swimtime="00:07:14.10" />
                    <SPLIT distance="725" swimtime="00:07:30.09" />
                    <SPLIT distance="750" swimtime="00:07:45.85" />
                    <SPLIT distance="775" swimtime="00:08:02.14" />
                    <SPLIT distance="800" swimtime="00:08:17.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154255" lastname="MILADINOV" firstname="Josif" gender="M" birthdate="2003-06-23">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.20" eventid="5" heat="6" lane="4">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="23" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="34" lane="4" heat="6" heatid="60005" swimtime="00:00:23.17" reactiontime="+64" points="827">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.76" />
                    <SPLIT distance="50" swimtime="00:00:23.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="25" lane="4" heat="1" heatid="10023" swimtime="00:00:54.06" reactiontime="+65" points="757">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.79" />
                    <SPLIT distance="50" swimtime="00:00:24.05" />
                    <SPLIT distance="75" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:00:54.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115408" lastname="GEORGIEVA" firstname="Gabriela" gender="F" birthdate="1997-06-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.94" eventid="2" heat="3" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.52" eventid="45" heat="2" lane="4">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="30" lane="2" heat="3" heatid="30002" swimtime="00:00:59.84" reactiontime="+61" points="771">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="75" swimtime="00:00:44.24" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="21" lane="4" heat="2" heatid="20045" swimtime="00:02:07.25" reactiontime="+61" points="816">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.49" />
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="75" swimtime="00:00:45.70" />
                    <SPLIT distance="100" swimtime="00:01:01.64" />
                    <SPLIT distance="125" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:01:34.00" />
                    <SPLIT distance="175" swimtime="00:01:50.59" />
                    <SPLIT distance="200" swimtime="00:02:07.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105114" lastname="PETKOVA" firstname="Diana" gender="F" birthdate="2000-06-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.05" eventid="13" heat="6" lane="4">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.98" eventid="40" heat="4" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.86" eventid="30" heat="7" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.58" eventid="22" heat="3" lane="6">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="31" lane="4" heat="6" heatid="60013" swimtime="00:00:54.58" reactiontime="+72" points="780">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="75" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:00:54.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="-1" lane="6" heat="4" heatid="40040" swimtime="00:00:30.61" status="DSQ" reactiontime="+71" />
                <RESULT eventid="30" place="23" lane="1" heat="7" heatid="70030" swimtime="00:00:24.96" reactiontime="+71" points="775">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                    <SPLIT distance="50" swimtime="00:00:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="15" lane="6" heat="3" heatid="30022" swimtime="00:01:00.08" reactiontime="+71" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.48" />
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                    <SPLIT distance="75" swimtime="00:00:45.20" />
                    <SPLIT distance="100" swimtime="00:01:00.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="11" lane="8" heat="2" heatid="20222" swimtime="00:00:59.45" reactiontime="+72" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                    <SPLIT distance="75" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Bulgaria">
              <RESULTS>
                <RESULT eventid="9" place="10" lane="1" heat="2" swimtime="00:03:12.15" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.78" />
                    <SPLIT distance="50" swimtime="00:00:22.55" />
                    <SPLIT distance="75" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:00:47.81" />
                    <SPLIT distance="125" swimtime="00:00:58.17" />
                    <SPLIT distance="150" swimtime="00:01:10.25" />
                    <SPLIT distance="175" swimtime="00:01:22.98" />
                    <SPLIT distance="200" swimtime="00:01:35.97" />
                    <SPLIT distance="225" swimtime="00:01:46.62" />
                    <SPLIT distance="250" swimtime="00:01:58.72" />
                    <SPLIT distance="275" swimtime="00:02:11.37" />
                    <SPLIT distance="300" swimtime="00:02:24.11" />
                    <SPLIT distance="325" swimtime="00:02:34.81" />
                    <SPLIT distance="350" swimtime="00:02:47.12" />
                    <SPLIT distance="375" swimtime="00:02:59.75" />
                    <SPLIT distance="400" swimtime="00:03:12.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202468" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="154255" reactiontime="+26" />
                    <RELAYPOSITION number="3" athleteid="105113" reactiontime="+4" />
                    <RELAYPOSITION number="4" athleteid="142443" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Bulgaria">
              <RESULTS>
                <RESULT eventid="48" place="14" lane="8" heat="2" swimtime="00:03:33.05" reactiontime="+52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="75" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:00:55.02" />
                    <SPLIT distance="125" swimtime="00:01:06.75" />
                    <SPLIT distance="150" swimtime="00:01:21.81" />
                    <SPLIT distance="175" swimtime="00:01:37.31" />
                    <SPLIT distance="200" swimtime="00:01:53.44" />
                    <SPLIT distance="225" swimtime="00:02:04.36" />
                    <SPLIT distance="250" swimtime="00:02:17.54" />
                    <SPLIT distance="275" swimtime="00:02:31.24" />
                    <SPLIT distance="300" swimtime="00:02:45.32" />
                    <SPLIT distance="325" swimtime="00:02:55.94" />
                    <SPLIT distance="350" swimtime="00:03:07.75" />
                    <SPLIT distance="375" swimtime="00:03:20.28" />
                    <SPLIT distance="400" swimtime="00:03:33.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="163143" reactiontime="+52" />
                    <RELAYPOSITION number="2" athleteid="213077" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="105113" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="202468" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Bulgaria">
              <RESULTS>
                <RESULT eventid="132" place="8" lane="7" heat="1" swimtime="00:06:59.12" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:24.09" />
                    <SPLIT distance="75" swimtime="00:00:37.11" />
                    <SPLIT distance="100" swimtime="00:00:50.52" />
                    <SPLIT distance="125" swimtime="00:01:03.71" />
                    <SPLIT distance="150" swimtime="00:01:17.26" />
                    <SPLIT distance="175" swimtime="00:01:30.97" />
                    <SPLIT distance="200" swimtime="00:01:44.31" />
                    <SPLIT distance="225" swimtime="00:01:54.88" />
                    <SPLIT distance="250" swimtime="00:02:07.78" />
                    <SPLIT distance="275" swimtime="00:02:20.87" />
                    <SPLIT distance="300" swimtime="00:02:34.43" />
                    <SPLIT distance="325" swimtime="00:02:47.36" />
                    <SPLIT distance="350" swimtime="00:03:00.90" />
                    <SPLIT distance="375" swimtime="00:03:14.69" />
                    <SPLIT distance="400" swimtime="00:03:28.24" />
                    <SPLIT distance="425" swimtime="00:03:39.13" />
                    <SPLIT distance="450" swimtime="00:03:51.99" />
                    <SPLIT distance="475" swimtime="00:04:05.47" />
                    <SPLIT distance="500" swimtime="00:04:18.99" />
                    <SPLIT distance="525" swimtime="00:04:32.59" />
                    <SPLIT distance="550" swimtime="00:04:46.08" />
                    <SPLIT distance="575" swimtime="00:04:59.55" />
                    <SPLIT distance="600" swimtime="00:05:12.69" />
                    <SPLIT distance="625" swimtime="00:05:24.10" />
                    <SPLIT distance="650" swimtime="00:05:37.08" />
                    <SPLIT distance="675" swimtime="00:05:50.20" />
                    <SPLIT distance="700" swimtime="00:06:03.58" />
                    <SPLIT distance="725" swimtime="00:06:16.95" />
                    <SPLIT distance="750" swimtime="00:06:30.64" />
                    <SPLIT distance="775" swimtime="00:06:45.04" />
                    <SPLIT distance="800" swimtime="00:06:59.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213076" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="142443" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="105113" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="149077" reactiontime="+3" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="6" lane="2" heat="2" swimtime="00:06:56.42" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.46" />
                    <SPLIT distance="50" swimtime="00:00:24.07" />
                    <SPLIT distance="75" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:00:50.07" />
                    <SPLIT distance="125" swimtime="00:01:03.28" />
                    <SPLIT distance="150" swimtime="00:01:16.72" />
                    <SPLIT distance="175" swimtime="00:01:30.44" />
                    <SPLIT distance="200" swimtime="00:01:43.76" />
                    <SPLIT distance="225" swimtime="00:01:54.80" />
                    <SPLIT distance="250" swimtime="00:02:07.80" />
                    <SPLIT distance="275" swimtime="00:02:21.24" />
                    <SPLIT distance="300" swimtime="00:02:34.76" />
                    <SPLIT distance="325" swimtime="00:02:47.66" />
                    <SPLIT distance="350" swimtime="00:03:00.68" />
                    <SPLIT distance="375" swimtime="00:03:14.19" />
                    <SPLIT distance="400" swimtime="00:03:27.44" />
                    <SPLIT distance="425" swimtime="00:03:38.44" />
                    <SPLIT distance="450" swimtime="00:03:51.01" />
                    <SPLIT distance="475" swimtime="00:04:03.90" />
                    <SPLIT distance="500" swimtime="00:04:17.33" />
                    <SPLIT distance="525" swimtime="00:04:30.68" />
                    <SPLIT distance="550" swimtime="00:04:44.08" />
                    <SPLIT distance="575" swimtime="00:04:57.78" />
                    <SPLIT distance="600" swimtime="00:05:10.99" />
                    <SPLIT distance="625" swimtime="00:05:22.50" />
                    <SPLIT distance="650" swimtime="00:05:35.43" />
                    <SPLIT distance="675" swimtime="00:05:48.68" />
                    <SPLIT distance="700" swimtime="00:06:02.02" />
                    <SPLIT distance="725" swimtime="00:06:15.43" />
                    <SPLIT distance="750" swimtime="00:06:29.04" />
                    <SPLIT distance="775" swimtime="00:06:42.81" />
                    <SPLIT distance="800" swimtime="00:06:56.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213076" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="142443" reactiontime="+37" />
                    <RELAYPOSITION number="3" athleteid="105113" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="149077" reactiontime="+4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Bulgaria">
              <RESULTS>
                <RESULT eventid="26" place="9" lane="1" heat="2" swimtime="00:01:26.58" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.15" />
                    <SPLIT distance="75" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:00:43.53" />
                    <SPLIT distance="125" swimtime="00:00:53.48" />
                    <SPLIT distance="150" swimtime="00:01:04.74" />
                    <SPLIT distance="175" swimtime="00:01:15.18" />
                    <SPLIT distance="200" swimtime="00:01:26.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154255" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="202468" reactiontime="+45" />
                    <RELAYPOSITION number="3" athleteid="142443" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="105113" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Bulgaria">
              <RESULTS>
                <RESULT eventid="11" place="13" lane="2" heat="3" swimtime="00:01:41.37" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="75" swimtime="00:00:39.30" />
                    <SPLIT distance="100" swimtime="00:00:53.80" />
                    <SPLIT distance="125" swimtime="00:01:04.10" />
                    <SPLIT distance="150" swimtime="00:01:16.87" />
                    <SPLIT distance="175" swimtime="00:01:28.57" />
                    <SPLIT distance="200" swimtime="00:01:41.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="115408" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="213077" reactiontime="0" />
                    <RELAYPOSITION number="3" athleteid="154255" reactiontime="+11" />
                    <RELAYPOSITION number="4" athleteid="105114" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Central African Rep" shortname="CAF" code="CAF" nation="CAF" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198080" lastname="TENGUE" firstname="Terence" gender="M" birthdate="2005-10-26">
              <ENTRIES>
                <ENTRY entrytime="00:00:34.27" eventid="31" heat="2" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="-1" lane="1" heat="2" heatid="20031" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Canada" shortname="CAN" code="CAN" nation="CAN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="124292" lastname="ACEVEDO" firstname="Javier" gender="M" birthdate="1998-01-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.71" eventid="3" heat="4" lane="5">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:01:49.74" eventid="46" heat="3" lane="5">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.80" eventid="7" heat="3" lane="6">
                  <MEETINFO date="2021-12-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:23.20" eventid="19" heat="4" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.38" eventid="23" heat="3" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="18" lane="5" heat="4" heatid="40003" swimtime="00:00:50.97" reactiontime="+56" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:24.81" />
                    <SPLIT distance="75" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:00:50.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="-1" lane="5" heat="3" heatid="30046" swimtime="00:01:50.50" status="DSQ" reactiontime="+57" />
                <RESULT eventid="7" place="17" lane="6" heat="3" heatid="30007" swimtime="00:01:54.96" reactiontime="+62" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.07" />
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                    <SPLIT distance="75" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:00:53.56" />
                    <SPLIT distance="125" swimtime="00:01:09.92" />
                    <SPLIT distance="150" swimtime="00:01:26.57" />
                    <SPLIT distance="175" swimtime="00:01:41.43" />
                    <SPLIT distance="200" swimtime="00:01:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="6" lane="3" heat="4" heatid="40019" swimtime="00:00:23.10" reactiontime="+56" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="8" lane="3" heat="1" heatid="10219" swimtime="00:00:23.05" reactiontime="+56" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="2" lane="3" heat="1" heatid="10123" swimtime="00:00:51.05" reactiontime="+60" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:23.43" />
                    <SPLIT distance="75" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:00:51.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="5" lane="4" heat="3" heatid="30023" swimtime="00:00:52.06" reactiontime="+59" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="75" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:00:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="3" lane="3" heat="2" heatid="20223" swimtime="00:00:51.46" reactiontime="+61" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.72" />
                    <SPLIT distance="50" swimtime="00:00:23.53" />
                    <SPLIT distance="75" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202149" lastname="DERGOUSOFF" firstname="James" gender="M" birthdate="1996-10-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.15" eventid="16" heat="4" lane="3">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.76" eventid="29" heat="2" lane="3">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:27.22" eventid="41" heat="6" lane="8">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="28" lane="3" heat="4" heatid="40016" swimtime="00:00:58.50" reactiontime="+69" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.75" />
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                    <SPLIT distance="75" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:00:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="13" lane="3" heat="2" heatid="20029" swimtime="00:02:06.17" reactiontime="+66" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="75" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:00.80" />
                    <SPLIT distance="125" swimtime="00:01:16.94" />
                    <SPLIT distance="150" swimtime="00:01:33.16" />
                    <SPLIT distance="175" swimtime="00:01:49.42" />
                    <SPLIT distance="200" swimtime="00:02:06.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="33" lane="8" heat="6" heatid="60041" swimtime="00:00:27.19" reactiontime="+68" points="772">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154453" lastname="KNOX" firstname="Finlay" gender="M" birthdate="2001-01-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.86" eventid="39" heat="4" lane="4">
                  <MEETINFO date="2022-04-06" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.32" eventid="7" heat="5" lane="3">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
                <ENTRY entrytime="00:04:07.09" eventid="37" heat="3" lane="7">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:51.70" eventid="23" heat="5" lane="3">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="-1" lane="4" heat="4" heatid="40039" swimtime="NT" status="DNS" />
                <RESULT eventid="107" place="3" lane="3" heat="1" heatid="10107" swimtime="00:01:51.04" reactiontime="+66" points="962">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.89" />
                    <SPLIT distance="50" swimtime="00:00:24.24" />
                    <SPLIT distance="75" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:00:52.32" />
                    <SPLIT distance="125" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:24.21" />
                    <SPLIT distance="175" swimtime="00:01:38.32" />
                    <SPLIT distance="200" swimtime="00:01:51.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="3" lane="3" heat="5" heatid="50007" swimtime="00:01:52.50" reactiontime="+67" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.84" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                    <SPLIT distance="75" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                    <SPLIT distance="125" swimtime="00:01:08.72" />
                    <SPLIT distance="150" swimtime="00:01:25.20" />
                    <SPLIT distance="175" swimtime="00:01:39.63" />
                    <SPLIT distance="200" swimtime="00:01:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="9" lane="7" heat="3" heatid="30037" swimtime="00:04:07.12" reactiontime="+67" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.11" />
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                    <SPLIT distance="75" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:00:54.65" />
                    <SPLIT distance="125" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:27.12" />
                    <SPLIT distance="175" swimtime="00:01:43.30" />
                    <SPLIT distance="200" swimtime="00:01:59.35" />
                    <SPLIT distance="225" swimtime="00:02:16.39" />
                    <SPLIT distance="250" swimtime="00:02:33.64" />
                    <SPLIT distance="275" swimtime="00:02:50.92" />
                    <SPLIT distance="300" swimtime="00:03:08.44" />
                    <SPLIT distance="325" swimtime="00:03:23.86" />
                    <SPLIT distance="350" swimtime="00:03:38.50" />
                    <SPLIT distance="375" swimtime="00:03:53.07" />
                    <SPLIT distance="400" swimtime="00:04:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="3" lane="7" heat="1" heatid="10123" swimtime="00:00:51.10" reactiontime="+66" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.42" />
                    <SPLIT distance="50" swimtime="00:00:23.09" />
                    <SPLIT distance="75" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:00:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="2" lane="3" heat="5" heatid="50023" swimtime="00:00:51.95" reactiontime="+70" points="853">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.71" />
                    <SPLIT distance="50" swimtime="00:00:23.58" />
                    <SPLIT distance="75" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:00:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="6" lane="4" heat="1" heatid="10223" swimtime="00:00:51.64" reactiontime="+66" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.55" />
                    <SPLIT distance="50" swimtime="00:00:23.33" />
                    <SPLIT distance="75" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214502" lastname="KHARUN" firstname="Ilya" gender="M" birthdate="2005-02-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.93" eventid="39" heat="7" lane="2">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.70" eventid="21" heat="4" lane="2">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:22.47" eventid="5" heat="8" lane="6">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="2" lane="2" heat="1" heatid="10139" swimtime="00:00:49.03" reactiontime="+66" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.65" />
                    <SPLIT distance="50" swimtime="00:00:23.11" />
                    <SPLIT distance="75" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:00:49.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="4" lane="2" heat="7" heatid="70039" swimtime="00:00:49.66" reactiontime="+67" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.29" />
                    <SPLIT distance="75" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:00:49.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="5" lane="5" heat="1" heatid="10239" swimtime="00:00:49.65" reactiontime="+69" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.72" />
                    <SPLIT distance="50" swimtime="00:00:23.16" />
                    <SPLIT distance="75" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:00:49.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="121" place="8" lane="1" heat="1" heatid="10121" swimtime="00:01:52.21" reactiontime="+67" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.07" />
                    <SPLIT distance="50" swimtime="00:00:24.98" />
                    <SPLIT distance="75" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:00:53.33" />
                    <SPLIT distance="125" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:22.31" />
                    <SPLIT distance="175" swimtime="00:01:37.26" />
                    <SPLIT distance="200" swimtime="00:01:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="7" lane="2" heat="4" heatid="40021" swimtime="00:01:50.86" reactiontime="+70" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.32" />
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                    <SPLIT distance="75" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:00:54.10" />
                    <SPLIT distance="125" swimtime="00:01:08.43" />
                    <SPLIT distance="150" swimtime="00:01:22.68" />
                    <SPLIT distance="175" swimtime="00:01:37.00" />
                    <SPLIT distance="200" swimtime="00:01:50.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="8" lane="6" heat="8" heatid="80005" swimtime="00:00:22.32" reactiontime="+68" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.42" />
                    <SPLIT distance="50" swimtime="00:00:22.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="8" lane="6" heat="1" heatid="10205" swimtime="00:00:22.28" reactiontime="+67" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.34" />
                    <SPLIT distance="50" swimtime="00:00:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="405" place="9" lane="4" heat="1" heatid="10405" swimtime="00:00:22.28" reactiontime="+63" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.26" />
                    <SPLIT distance="50" swimtime="00:00:22.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118562" lastname="KISIL" firstname="Yuri" gender="M" birthdate="1995-09-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.09" eventid="14" heat="11" lane="8">
                  <MEETINFO date="2021-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:21.37" eventid="31" heat="9" lane="1">
                  <MEETINFO date="2021-09-10" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="28" lane="8" heat="11" heatid="110014" swimtime="00:00:47.40" reactiontime="+69" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.83" />
                    <SPLIT distance="50" swimtime="00:00:22.83" />
                    <SPLIT distance="75" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="65" lane="1" heat="9" heatid="90031" swimtime="00:00:25.14" reactiontime="+67" points="515">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:25.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149353" lastname="GAZIEV" firstname="Ruslan" gender="M" birthdate="1999-08-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.41" eventid="14" heat="7" lane="7">
                  <MEETINFO date="2022-04-08" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.44" eventid="44" heat="2" lane="5">
                  <MEETINFO date="2022-04-07" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="25" lane="7" heat="7" heatid="70014" swimtime="00:00:47.30" reactiontime="+65" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.44" />
                    <SPLIT distance="75" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="23" lane="5" heat="2" heatid="20044" swimtime="00:01:44.97" reactiontime="+66" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:24.69" />
                    <SPLIT distance="75" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:00:51.45" />
                    <SPLIT distance="125" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:18.24" />
                    <SPLIT distance="175" swimtime="00:01:31.97" />
                    <SPLIT distance="200" swimtime="00:01:44.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129652" lastname="MASSE" firstname="Kylie" gender="F" birthdate="1996-01-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.22" eventid="2" heat="5" lane="4">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.45" eventid="45" heat="5" lane="5">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:25.62" eventid="18" heat="6" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="6" lane="2" heat="1" heatid="10102" swimtime="00:00:56.18" reactiontime="+58" points="932">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.21" />
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="75" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:00:56.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="10" lane="4" heat="5" heatid="50002" swimtime="00:00:57.01" reactiontime="+57" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="75" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:00:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="5" lane="7" heat="2" heatid="20202" swimtime="00:00:56.13" reactiontime="+58" points="935">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                    <SPLIT distance="75" swimtime="00:00:41.53" />
                    <SPLIT distance="100" swimtime="00:00:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="3" lane="3" heat="1" heatid="10145" swimtime="00:02:01.26" reactiontime="+60" points="943">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="75" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                    <SPLIT distance="125" swimtime="00:01:14.85" />
                    <SPLIT distance="150" swimtime="00:01:30.32" />
                    <SPLIT distance="175" swimtime="00:01:45.97" />
                    <SPLIT distance="200" swimtime="00:02:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="3" lane="5" heat="5" heatid="50045" swimtime="00:02:02.54" reactiontime="+55" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="75" swimtime="00:00:44.56" />
                    <SPLIT distance="100" swimtime="00:01:00.14" />
                    <SPLIT distance="125" swimtime="00:01:15.63" />
                    <SPLIT distance="150" swimtime="00:01:31.43" />
                    <SPLIT distance="175" swimtime="00:01:47.32" />
                    <SPLIT distance="200" swimtime="00:02:02.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="4" lane="6" heat="1" heatid="10118" swimtime="00:00:25.81" reactiontime="+58" points="938">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="2" lane="4" heat="6" heatid="60018" swimtime="00:00:25.94" reactiontime="+56" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.83" />
                    <SPLIT distance="50" swimtime="00:00:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="4" lane="4" heat="1" heatid="10218" swimtime="00:00:25.97" reactiontime="+57" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156529" lastname="WILM" firstname="Ingrid" gender="F" birthdate="1998-06-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.61" eventid="2" heat="6" lane="5">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.26" eventid="45" heat="5" lane="3">
                  <MEETINFO date="2021-09-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="3" lane="5" heat="1" heatid="10102" swimtime="00:00:55.74" reactiontime="+65" points="954">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="75" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:00:55.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="2" lane="5" heat="6" heatid="60002" swimtime="00:00:56.15" reactiontime="+64" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="75" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:00:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="2" lane="4" heat="1" heatid="10202" swimtime="00:00:55.92" reactiontime="+63" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="75" swimtime="00:00:41.47" />
                    <SPLIT distance="100" swimtime="00:00:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="4" lane="8" heat="1" heatid="10145" swimtime="00:02:01.78" reactiontime="+65" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="75" swimtime="00:00:44.83" />
                    <SPLIT distance="100" swimtime="00:01:00.79" />
                    <SPLIT distance="125" swimtime="00:01:16.18" />
                    <SPLIT distance="150" swimtime="00:01:31.37" />
                    <SPLIT distance="175" swimtime="00:01:46.82" />
                    <SPLIT distance="200" swimtime="00:02:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="8" lane="3" heat="5" heatid="50045" swimtime="00:02:03.57" reactiontime="+62" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                    <SPLIT distance="75" swimtime="00:00:45.57" />
                    <SPLIT distance="100" swimtime="00:01:01.52" />
                    <SPLIT distance="125" swimtime="00:01:17.42" />
                    <SPLIT distance="150" swimtime="00:01:32.96" />
                    <SPLIT distance="175" swimtime="00:01:48.52" />
                    <SPLIT distance="200" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118565" lastname="NICOL" firstname="Rachel" gender="F" birthdate="1993-02-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.01" eventid="15" heat="4" lane="6">
                  <MEETINFO date="2021-11-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:30.84" eventid="40" heat="4" lane="5">
                  <MEETINFO date="2021-11-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="24" lane="6" heat="4" heatid="40015" swimtime="00:01:05.91" reactiontime="+66" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.49" />
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="75" swimtime="00:00:48.47" />
                    <SPLIT distance="100" swimtime="00:01:05.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="20" lane="5" heat="4" heatid="40040" swimtime="00:00:30.43" reactiontime="+63" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.19" />
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118566" lastname="PICKREM" firstname="Sydney" gender="F" birthdate="1997-05-21">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.38" eventid="15" heat="7" lane="1">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.71" eventid="28" heat="3" lane="5">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.29" eventid="6" heat="4" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:04:26.66" eventid="36" heat="3" lane="4">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:00:58.40" eventid="22" heat="3" lane="5">
                  <MEETINFO date="2021-09-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="10" lane="1" heat="7" heatid="70015" swimtime="00:01:04.73" reactiontime="+69" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.11" />
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="75" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:04.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="12" lane="2" heat="1" heatid="10215" swimtime="00:01:05.08" reactiontime="+67" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="75" swimtime="00:00:47.82" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="128" place="6" lane="6" heat="1" heatid="10128" swimtime="00:02:19.35" reactiontime="+73" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.49" />
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="75" swimtime="00:00:49.29" />
                    <SPLIT distance="100" swimtime="00:01:06.92" />
                    <SPLIT distance="125" swimtime="00:01:24.85" />
                    <SPLIT distance="150" swimtime="00:01:42.95" />
                    <SPLIT distance="175" swimtime="00:02:01.10" />
                    <SPLIT distance="200" swimtime="00:02:19.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="4" lane="5" heat="3" heatid="30028" swimtime="00:02:19.57" reactiontime="+73" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="75" swimtime="00:00:49.72" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="125" swimtime="00:01:25.58" />
                    <SPLIT distance="150" swimtime="00:01:43.61" />
                    <SPLIT distance="175" swimtime="00:02:01.62" />
                    <SPLIT distance="200" swimtime="00:02:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106" place="5" lane="7" heat="1" heatid="10106" swimtime="00:02:05.22" reactiontime="+75" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="75" swimtime="00:00:43.81" />
                    <SPLIT distance="100" swimtime="00:00:59.11" />
                    <SPLIT distance="125" swimtime="00:01:16.75" />
                    <SPLIT distance="150" swimtime="00:01:34.98" />
                    <SPLIT distance="175" swimtime="00:01:50.67" />
                    <SPLIT distance="200" swimtime="00:02:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="6" lane="4" heat="4" heatid="40006" swimtime="00:02:07.15" reactiontime="+67" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                    <SPLIT distance="75" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:00.12" />
                    <SPLIT distance="125" swimtime="00:01:18.43" />
                    <SPLIT distance="150" swimtime="00:01:36.66" />
                    <SPLIT distance="175" swimtime="00:01:52.51" />
                    <SPLIT distance="200" swimtime="00:02:07.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="-1" lane="4" heat="3" heatid="30036" swimtime="NT" status="DNS" />
                <RESULT eventid="122" place="4" lane="3" heat="1" heatid="10122" swimtime="00:00:58.26" reactiontime="+67" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                    <SPLIT distance="75" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:00:58.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="10" lane="5" heat="3" heatid="30022" swimtime="00:00:59.49" reactiontime="+70" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.61" />
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="75" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="3" lane="7" heat="2" heatid="20222" swimtime="00:00:58.54" reactiontime="+71" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="75" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:00:58.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101207" lastname="SAVARD" firstname="Katerine" gender="F" birthdate="1993-05-26">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.23" eventid="38" heat="4" lane="7">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.15" eventid="13" heat="9" lane="7">
                  <MEETINFO date="2021-12-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.64" eventid="20" heat="2" lane="3">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:00:26.14" eventid="4" heat="6" lane="7">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="138" place="8" lane="1" heat="1" heatid="10138" swimtime="00:00:56.87" reactiontime="+63" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.09" />
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                    <SPLIT distance="75" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:00:56.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="8" lane="7" heat="4" heatid="40038" swimtime="00:00:56.86" reactiontime="+65" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="75" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:00:56.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="8" lane="6" heat="1" heatid="10238" swimtime="00:00:56.44" reactiontime="+63" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.03" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="75" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:00:56.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="19" lane="7" heat="9" heatid="90013" swimtime="00:00:53.59" reactiontime="+62" points="824">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                    <SPLIT distance="50" swimtime="00:00:25.88" />
                    <SPLIT distance="75" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:00:53.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="14" lane="3" heat="2" heatid="20020" swimtime="00:02:08.51" reactiontime="+65" points="806">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.96" />
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="75" swimtime="00:00:44.77" />
                    <SPLIT distance="100" swimtime="00:01:01.00" />
                    <SPLIT distance="125" swimtime="00:01:17.03" />
                    <SPLIT distance="150" swimtime="00:01:33.40" />
                    <SPLIT distance="175" swimtime="00:01:50.19" />
                    <SPLIT distance="200" swimtime="00:02:08.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="13" lane="7" heat="6" heatid="60004" swimtime="00:00:25.50" reactiontime="+62" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="16" lane="1" heat="2" heatid="20204" swimtime="00:00:25.81" reactiontime="+64" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124174" lastname="MACNEIL" firstname="Margaret" gender="F" birthdate="2000-02-26">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.78" eventid="38" heat="4" lane="4">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:25.27" eventid="18" heat="7" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.75" eventid="4" heat="5" lane="4">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="138" place="1" lane="3" heat="1" heatid="10138" swimtime="00:00:54.05" reactiontime="+62" points="1030">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.69" />
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                    <SPLIT distance="75" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="4" lane="4" heat="4" heatid="40038" swimtime="00:00:56.53" reactiontime="+57" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                    <SPLIT distance="75" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:00:56.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="3" lane="5" heat="1" heatid="10238" swimtime="00:00:55.83" reactiontime="+66" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="75" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:00:55.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="1" lane="5" heat="1" heatid="10118" swimtime="00:00:25.25" reactiontime="+56" points="1002">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="7" lane="4" heat="7" heatid="70018" swimtime="00:00:26.09" reactiontime="+58" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="2" lane="6" heat="1" heatid="10218" swimtime="00:00:25.64" reactiontime="+58" points="957">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="104" place="1" lane="4" heat="1" heatid="10104" swimtime="00:00:24.64" reactiontime="+64" points="968">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="5" lane="4" heat="5" heatid="50004" swimtime="00:00:25.13" reactiontime="+67" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="1" lane="3" heat="2" heatid="20204" swimtime="00:00:24.78" reactiontime="+65" points="952">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                    <SPLIT distance="50" swimtime="00:00:24.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124058" lastname="RUCK" firstname="Taylor" gender="F" birthdate="2000-05-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.99" eventid="13" heat="7" lane="8">
                  <MEETINFO date="2022-04-08" />
                </ENTRY>
                <ENTRY entrytime="00:01:56.80" eventid="43" heat="5" lane="7">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="6" lane="8" heat="1" heatid="10113" swimtime="00:00:52.08" reactiontime="+68" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="75" swimtime="00:00:38.34" />
                    <SPLIT distance="100" swimtime="00:00:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="8" lane="8" heat="7" heatid="70013" swimtime="00:00:52.56" reactiontime="+70" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:25.15" />
                    <SPLIT distance="75" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:00:52.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="8" lane="6" heat="1" heatid="10213" swimtime="00:00:52.27" reactiontime="+69" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:25.06" />
                    <SPLIT distance="75" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:00:52.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="143" place="7" lane="1" heat="1" heatid="10143" swimtime="00:01:52.88" reactiontime="+66" points="933">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.27" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:54.74" />
                    <SPLIT distance="125" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:23.79" />
                    <SPLIT distance="175" swimtime="00:01:38.45" />
                    <SPLIT distance="200" swimtime="00:01:52.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="7" lane="7" heat="5" heatid="50043" swimtime="00:01:54.15" reactiontime="+70" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="75" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:00:55.70" />
                    <SPLIT distance="125" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:24.72" />
                    <SPLIT distance="175" swimtime="00:01:39.54" />
                    <SPLIT distance="200" swimtime="00:01:54.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129690" lastname="WOG" firstname="Kelsey Lauren" gender="F" birthdate="1998-09-19">
              <ENTRIES>
                <ENTRY entrytime="00:02:20.59" eventid="28" heat="5" lane="6">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="10" lane="6" heat="5" heatid="50028" swimtime="00:02:20.57" reactiontime="+66" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="75" swimtime="00:00:49.62" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="125" swimtime="00:01:25.75" />
                    <SPLIT distance="150" swimtime="00:01:43.82" />
                    <SPLIT distance="175" swimtime="00:02:02.06" />
                    <SPLIT distance="200" swimtime="00:02:20.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124394" lastname="SMITH" firstname="Rebecca" gender="F" birthdate="2000-03-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.24" eventid="43" heat="5" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="143" place="2" lane="2" heat="1" heatid="10143" swimtime="00:01:52.24" reactiontime="+71" points="949">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="75" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:00:54.41" />
                    <SPLIT distance="125" swimtime="00:01:08.78" />
                    <SPLIT distance="150" swimtime="00:01:23.19" />
                    <SPLIT distance="175" swimtime="00:01:37.82" />
                    <SPLIT distance="200" swimtime="00:01:52.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="5" lane="5" heat="5" heatid="50043" swimtime="00:01:53.85" reactiontime="+71" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                    <SPLIT distance="75" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:00:55.92" />
                    <SPLIT distance="125" swimtime="00:01:10.39" />
                    <SPLIT distance="150" swimtime="00:01:25.03" />
                    <SPLIT distance="175" swimtime="00:01:39.71" />
                    <SPLIT distance="200" swimtime="00:01:53.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124399" lastname="HARVEY" firstname="Mary-Sophie" gender="F" birthdate="1999-08-11">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.15" eventid="6" heat="4" lane="5">
                  <MEETINFO date="2021-09-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:00:58.24" eventid="22" heat="4" lane="5">
                  <MEETINFO date="2021-11-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="9" lane="5" heat="4" heatid="40006" swimtime="00:02:07.41" reactiontime="+67" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="75" swimtime="00:00:44.70" />
                    <SPLIT distance="100" swimtime="00:01:00.60" />
                    <SPLIT distance="125" swimtime="00:01:18.90" />
                    <SPLIT distance="150" swimtime="00:01:37.56" />
                    <SPLIT distance="175" swimtime="00:01:53.25" />
                    <SPLIT distance="200" swimtime="00:02:07.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="8" lane="1" heat="1" heatid="10122" swimtime="00:00:59.11" reactiontime="+67" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                    <SPLIT distance="75" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:00:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="4" lane="5" heat="4" heatid="40022" swimtime="00:00:58.93" reactiontime="+66" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.27" />
                    <SPLIT distance="50" swimtime="00:00:26.63" />
                    <SPLIT distance="75" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:00:58.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="7" lane="5" heat="1" heatid="10222" swimtime="00:00:59.13" reactiontime="+67" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                    <SPLIT distance="75" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124173" lastname="CIEPLUCHA" firstname="Tessa" gender="F" birthdate="1998-09-24">
              <ENTRIES>
                <ENTRY entrytime="00:04:25.55" eventid="36" heat="4" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="136" place="-1" lane="1" heat="1" heatid="10136" swimtime="00:04:34.79" status="DSQ" reactiontime="+77" />
                <RESULT eventid="36" place="7" lane="4" heat="4" heatid="40036" swimtime="00:04:33.58" reactiontime="+74" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="75" swimtime="00:00:45.51" />
                    <SPLIT distance="100" swimtime="00:01:02.31" />
                    <SPLIT distance="125" swimtime="00:01:20.53" />
                    <SPLIT distance="150" swimtime="00:01:37.99" />
                    <SPLIT distance="175" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:12.65" />
                    <SPLIT distance="225" swimtime="00:02:31.73" />
                    <SPLIT distance="250" swimtime="00:02:50.82" />
                    <SPLIT distance="275" swimtime="00:03:10.47" />
                    <SPLIT distance="300" swimtime="00:03:30.15" />
                    <SPLIT distance="325" swimtime="00:03:46.78" />
                    <SPLIT distance="350" swimtime="00:04:02.59" />
                    <SPLIT distance="375" swimtime="00:04:18.41" />
                    <SPLIT distance="400" swimtime="00:04:33.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Canada">
              <RESULTS>
                <RESULT eventid="109" place="5" lane="1" heat="1" swimtime="00:03:07.10" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.43" />
                    <SPLIT distance="75" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:00:47.08" />
                    <SPLIT distance="125" swimtime="00:00:57.40" />
                    <SPLIT distance="150" swimtime="00:01:09.32" />
                    <SPLIT distance="175" swimtime="00:01:21.52" />
                    <SPLIT distance="200" swimtime="00:01:33.49" />
                    <SPLIT distance="225" swimtime="00:01:43.62" />
                    <SPLIT distance="250" swimtime="00:01:55.38" />
                    <SPLIT distance="275" swimtime="00:02:07.58" />
                    <SPLIT distance="300" swimtime="00:02:19.67" />
                    <SPLIT distance="325" swimtime="00:02:29.75" />
                    <SPLIT distance="350" swimtime="00:02:41.95" />
                    <SPLIT distance="375" swimtime="00:02:54.75" />
                    <SPLIT distance="400" swimtime="00:03:07.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="149353" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="118562" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="124292" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="214502" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="7" lane="6" heat="2" swimtime="00:03:08.80" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.67" />
                    <SPLIT distance="50" swimtime="00:00:22.55" />
                    <SPLIT distance="75" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:00:47.32" />
                    <SPLIT distance="125" swimtime="00:00:57.49" />
                    <SPLIT distance="150" swimtime="00:01:09.53" />
                    <SPLIT distance="175" swimtime="00:01:22.26" />
                    <SPLIT distance="200" swimtime="00:01:34.66" />
                    <SPLIT distance="225" swimtime="00:01:44.95" />
                    <SPLIT distance="250" swimtime="00:01:56.91" />
                    <SPLIT distance="275" swimtime="00:02:09.04" />
                    <SPLIT distance="300" swimtime="00:02:21.23" />
                    <SPLIT distance="325" swimtime="00:02:31.71" />
                    <SPLIT distance="350" swimtime="00:02:43.97" />
                    <SPLIT distance="375" swimtime="00:02:56.61" />
                    <SPLIT distance="400" swimtime="00:03:08.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="149353" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="214502" reactiontime="+8" />
                    <RELAYPOSITION number="3" athleteid="118562" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="154453" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Canada">
              <RESULTS>
                <RESULT eventid="148" place="6" lane="7" heat="1" swimtime="00:03:23.44" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.69" />
                    <SPLIT distance="50" swimtime="00:00:24.17" />
                    <SPLIT distance="75" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:00:50.46" />
                    <SPLIT distance="125" swimtime="00:01:01.90" />
                    <SPLIT distance="150" swimtime="00:01:16.69" />
                    <SPLIT distance="175" swimtime="00:01:31.83" />
                    <SPLIT distance="200" swimtime="00:01:47.67" />
                    <SPLIT distance="225" swimtime="00:01:57.83" />
                    <SPLIT distance="250" swimtime="00:02:10.74" />
                    <SPLIT distance="275" swimtime="00:02:23.87" />
                    <SPLIT distance="300" swimtime="00:02:37.21" />
                    <SPLIT distance="325" swimtime="00:02:47.22" />
                    <SPLIT distance="350" swimtime="00:02:59.02" />
                    <SPLIT distance="375" swimtime="00:03:11.27" />
                    <SPLIT distance="400" swimtime="00:03:23.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154453" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="124292" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="214502" reactiontime="+16" />
                    <RELAYPOSITION number="4" athleteid="149353" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="6" lane="7" heat="3" swimtime="00:03:25.33" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:24.32" />
                    <SPLIT distance="75" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:00:50.40" />
                    <SPLIT distance="125" swimtime="00:01:02.88" />
                    <SPLIT distance="150" swimtime="00:01:17.60" />
                    <SPLIT distance="175" swimtime="00:01:32.66" />
                    <SPLIT distance="200" swimtime="00:01:48.78" />
                    <SPLIT distance="225" swimtime="00:01:58.84" />
                    <SPLIT distance="250" swimtime="00:02:11.64" />
                    <SPLIT distance="275" swimtime="00:02:24.94" />
                    <SPLIT distance="300" swimtime="00:02:38.54" />
                    <SPLIT distance="325" swimtime="00:02:48.88" />
                    <SPLIT distance="350" swimtime="00:03:00.74" />
                    <SPLIT distance="375" swimtime="00:03:13.00" />
                    <SPLIT distance="400" swimtime="00:03:25.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154453" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="202149" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="214502" reactiontime="+6" />
                    <RELAYPOSITION number="4" athleteid="118562" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Canada">
              <RESULTS>
                <RESULT eventid="132" place="7" lane="8" heat="1" swimtime="00:06:56.02" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.98" />
                    <SPLIT distance="50" swimtime="00:00:23.85" />
                    <SPLIT distance="75" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:00:50.67" />
                    <SPLIT distance="125" swimtime="00:01:03.95" />
                    <SPLIT distance="150" swimtime="00:01:17.48" />
                    <SPLIT distance="175" swimtime="00:01:30.94" />
                    <SPLIT distance="200" swimtime="00:01:43.96" />
                    <SPLIT distance="225" swimtime="00:01:54.71" />
                    <SPLIT distance="250" swimtime="00:02:07.76" />
                    <SPLIT distance="275" swimtime="00:02:21.08" />
                    <SPLIT distance="300" swimtime="00:02:34.65" />
                    <SPLIT distance="325" swimtime="00:02:48.01" />
                    <SPLIT distance="350" swimtime="00:03:01.42" />
                    <SPLIT distance="375" swimtime="00:03:14.95" />
                    <SPLIT distance="400" swimtime="00:03:28.28" />
                    <SPLIT distance="425" swimtime="00:03:38.80" />
                    <SPLIT distance="450" swimtime="00:03:52.08" />
                    <SPLIT distance="475" swimtime="00:04:05.68" />
                    <SPLIT distance="500" swimtime="00:04:19.31" />
                    <SPLIT distance="525" swimtime="00:04:33.01" />
                    <SPLIT distance="550" swimtime="00:04:46.79" />
                    <SPLIT distance="575" swimtime="00:05:00.49" />
                    <SPLIT distance="600" swimtime="00:05:13.79" />
                    <SPLIT distance="625" swimtime="00:05:24.09" />
                    <SPLIT distance="650" swimtime="00:05:36.47" />
                    <SPLIT distance="675" swimtime="00:05:49.05" />
                    <SPLIT distance="700" swimtime="00:06:02.12" />
                    <SPLIT distance="725" swimtime="00:06:15.33" />
                    <SPLIT distance="750" swimtime="00:06:28.68" />
                    <SPLIT distance="775" swimtime="00:06:42.47" />
                    <SPLIT distance="800" swimtime="00:06:56.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154453" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="149353" reactiontime="+35" />
                    <RELAYPOSITION number="3" athleteid="214502" reactiontime="+9" />
                    <RELAYPOSITION number="4" athleteid="124292" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="8" lane="6" heat="1" swimtime="00:07:00.85" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:24.57" />
                    <SPLIT distance="75" swimtime="00:00:37.90" />
                    <SPLIT distance="100" swimtime="00:00:51.13" />
                    <SPLIT distance="125" swimtime="00:01:04.60" />
                    <SPLIT distance="150" swimtime="00:01:18.04" />
                    <SPLIT distance="175" swimtime="00:01:31.67" />
                    <SPLIT distance="200" swimtime="00:01:44.73" />
                    <SPLIT distance="225" swimtime="00:01:55.61" />
                    <SPLIT distance="250" swimtime="00:02:08.83" />
                    <SPLIT distance="275" swimtime="00:02:22.48" />
                    <SPLIT distance="300" swimtime="00:02:36.06" />
                    <SPLIT distance="325" swimtime="00:02:49.88" />
                    <SPLIT distance="350" swimtime="00:03:03.52" />
                    <SPLIT distance="375" swimtime="00:03:17.29" />
                    <SPLIT distance="400" swimtime="00:03:30.16" />
                    <SPLIT distance="425" swimtime="00:03:41.30" />
                    <SPLIT distance="450" swimtime="00:03:54.70" />
                    <SPLIT distance="475" swimtime="00:04:08.24" />
                    <SPLIT distance="500" swimtime="00:04:21.89" />
                    <SPLIT distance="525" swimtime="00:04:35.45" />
                    <SPLIT distance="550" swimtime="00:04:49.18" />
                    <SPLIT distance="575" swimtime="00:05:02.84" />
                    <SPLIT distance="600" swimtime="00:05:16.18" />
                    <SPLIT distance="625" swimtime="00:05:26.84" />
                    <SPLIT distance="650" swimtime="00:05:39.59" />
                    <SPLIT distance="675" swimtime="00:05:52.74" />
                    <SPLIT distance="700" swimtime="00:06:06.11" />
                    <SPLIT distance="725" swimtime="00:06:19.71" />
                    <SPLIT distance="750" swimtime="00:06:33.49" />
                    <SPLIT distance="775" swimtime="00:06:47.47" />
                    <SPLIT distance="800" swimtime="00:07:00.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="149353" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="214502" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="118562" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="154453" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Canada">
              <RESULTS>
                <RESULT eventid="27" place="-1" lane="4" heat="4" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Canada">
              <RESULTS>
                <RESULT eventid="108" place="3" lane="3" heat="1" swimtime="00:03:28.06" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.08" />
                    <SPLIT distance="50" swimtime="00:00:25.32" />
                    <SPLIT distance="75" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:00:52.68" />
                    <SPLIT distance="125" swimtime="00:01:04.10" />
                    <SPLIT distance="150" swimtime="00:01:17.02" />
                    <SPLIT distance="175" swimtime="00:01:30.52" />
                    <SPLIT distance="200" swimtime="00:01:44.17" />
                    <SPLIT distance="225" swimtime="00:01:55.47" />
                    <SPLIT distance="250" swimtime="00:02:08.48" />
                    <SPLIT distance="275" swimtime="00:02:21.87" />
                    <SPLIT distance="300" swimtime="00:02:35.28" />
                    <SPLIT distance="325" swimtime="00:02:47.20" />
                    <SPLIT distance="350" swimtime="00:03:00.15" />
                    <SPLIT distance="375" swimtime="00:03:13.96" />
                    <SPLIT distance="400" swimtime="00:03:28.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124394" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="124058" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="124174" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="101207" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="3" lane="4" heat="2" swimtime="00:03:30.69" reactiontime="+71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.19" />
                    <SPLIT distance="50" swimtime="00:00:25.47" />
                    <SPLIT distance="75" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:00:52.75" />
                    <SPLIT distance="125" swimtime="00:01:04.80" />
                    <SPLIT distance="150" swimtime="00:01:18.15" />
                    <SPLIT distance="175" swimtime="00:01:31.85" />
                    <SPLIT distance="200" swimtime="00:01:45.65" />
                    <SPLIT distance="225" swimtime="00:01:57.79" />
                    <SPLIT distance="250" swimtime="00:02:11.16" />
                    <SPLIT distance="275" swimtime="00:02:24.99" />
                    <SPLIT distance="300" swimtime="00:02:38.78" />
                    <SPLIT distance="325" swimtime="00:02:50.22" />
                    <SPLIT distance="350" swimtime="00:03:03.41" />
                    <SPLIT distance="375" swimtime="00:03:17.13" />
                    <SPLIT distance="400" swimtime="00:03:30.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124394" reactiontime="+71" />
                    <RELAYPOSITION number="2" athleteid="101207" reactiontime="+45" />
                    <RELAYPOSITION number="3" athleteid="124399" reactiontime="+48" />
                    <RELAYPOSITION number="4" athleteid="124058" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Canada">
              <RESULTS>
                <RESULT eventid="147" place="3" lane="3" heat="1" swimtime="00:03:46.22" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                    <SPLIT distance="75" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:00:55.36" />
                    <SPLIT distance="125" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:25.58" />
                    <SPLIT distance="175" swimtime="00:01:42.54" />
                    <SPLIT distance="200" swimtime="00:01:59.78" />
                    <SPLIT distance="225" swimtime="00:02:10.98" />
                    <SPLIT distance="250" swimtime="00:02:24.87" />
                    <SPLIT distance="275" swimtime="00:02:39.37" />
                    <SPLIT distance="300" swimtime="00:02:54.37" />
                    <SPLIT distance="325" swimtime="00:03:05.69" />
                    <SPLIT distance="350" swimtime="00:03:18.71" />
                    <SPLIT distance="375" swimtime="00:03:32.28" />
                    <SPLIT distance="400" swimtime="00:03:46.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156529" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="118566" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="124174" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="124058" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="3" lane="4" heat="1" swimtime="00:03:51.40" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                    <SPLIT distance="75" swimtime="00:00:41.76" />
                    <SPLIT distance="100" swimtime="00:00:56.41" />
                    <SPLIT distance="125" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:26.93" />
                    <SPLIT distance="175" swimtime="00:01:44.13" />
                    <SPLIT distance="200" swimtime="00:02:01.85" />
                    <SPLIT distance="225" swimtime="00:02:13.84" />
                    <SPLIT distance="250" swimtime="00:02:28.24" />
                    <SPLIT distance="275" swimtime="00:02:43.34" />
                    <SPLIT distance="300" swimtime="00:02:59.06" />
                    <SPLIT distance="325" swimtime="00:03:10.87" />
                    <SPLIT distance="350" swimtime="00:03:24.24" />
                    <SPLIT distance="375" swimtime="00:03:37.89" />
                    <SPLIT distance="400" swimtime="00:03:51.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129652" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="118565" reactiontime="+36" />
                    <RELAYPOSITION number="3" athleteid="101207" reactiontime="+42" />
                    <RELAYPOSITION number="4" athleteid="124394" reactiontime="+41" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Canada">
              <RESULTS>
                <RESULT eventid="117" place="2" lane="2" heat="1" swimtime="00:07:34.47" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                    <SPLIT distance="75" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:00:54.41" />
                    <SPLIT distance="125" swimtime="00:01:08.75" />
                    <SPLIT distance="150" swimtime="00:01:23.28" />
                    <SPLIT distance="175" swimtime="00:01:37.81" />
                    <SPLIT distance="200" swimtime="00:01:52.15" />
                    <SPLIT distance="225" swimtime="00:02:04.46" />
                    <SPLIT distance="250" swimtime="00:02:18.34" />
                    <SPLIT distance="275" swimtime="00:02:32.81" />
                    <SPLIT distance="300" swimtime="00:02:47.48" />
                    <SPLIT distance="325" swimtime="00:03:02.15" />
                    <SPLIT distance="350" swimtime="00:03:17.04" />
                    <SPLIT distance="375" swimtime="00:03:32.08" />
                    <SPLIT distance="400" swimtime="00:03:46.93" />
                    <SPLIT distance="425" swimtime="00:03:59.05" />
                    <SPLIT distance="450" swimtime="00:04:12.89" />
                    <SPLIT distance="475" swimtime="00:04:27.00" />
                    <SPLIT distance="500" swimtime="00:04:41.61" />
                    <SPLIT distance="525" swimtime="00:04:56.34" />
                    <SPLIT distance="550" swimtime="00:05:11.36" />
                    <SPLIT distance="575" swimtime="00:05:26.66" />
                    <SPLIT distance="600" swimtime="00:05:41.74" />
                    <SPLIT distance="625" swimtime="00:05:53.49" />
                    <SPLIT distance="650" swimtime="00:06:07.09" />
                    <SPLIT distance="675" swimtime="00:06:21.11" />
                    <SPLIT distance="700" swimtime="00:06:35.48" />
                    <SPLIT distance="725" swimtime="00:06:49.80" />
                    <SPLIT distance="750" swimtime="00:07:04.43" />
                    <SPLIT distance="775" swimtime="00:07:19.42" />
                    <SPLIT distance="800" swimtime="00:07:34.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124394" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="101207" reactiontime="+45" />
                    <RELAYPOSITION number="3" athleteid="124399" reactiontime="+52" />
                    <RELAYPOSITION number="4" athleteid="124058" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="5" lane="4" heat="2" swimtime="00:07:46.70" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.83" />
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                    <SPLIT distance="75" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:00:56.70" />
                    <SPLIT distance="125" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:26.33" />
                    <SPLIT distance="175" swimtime="00:01:41.10" />
                    <SPLIT distance="200" swimtime="00:01:55.58" />
                    <SPLIT distance="225" swimtime="00:02:08.51" />
                    <SPLIT distance="250" swimtime="00:02:23.06" />
                    <SPLIT distance="275" swimtime="00:02:37.85" />
                    <SPLIT distance="300" swimtime="00:02:52.82" />
                    <SPLIT distance="325" swimtime="00:03:07.81" />
                    <SPLIT distance="350" swimtime="00:03:22.89" />
                    <SPLIT distance="375" swimtime="00:03:37.94" />
                    <SPLIT distance="400" swimtime="00:03:52.65" />
                    <SPLIT distance="425" swimtime="00:04:05.44" />
                    <SPLIT distance="450" swimtime="00:04:19.94" />
                    <SPLIT distance="475" swimtime="00:04:34.62" />
                    <SPLIT distance="500" swimtime="00:04:49.50" />
                    <SPLIT distance="525" swimtime="00:05:04.15" />
                    <SPLIT distance="550" swimtime="00:05:19.04" />
                    <SPLIT distance="575" swimtime="00:05:34.01" />
                    <SPLIT distance="600" swimtime="00:05:48.83" />
                    <SPLIT distance="625" swimtime="00:06:01.77" />
                    <SPLIT distance="650" swimtime="00:06:16.15" />
                    <SPLIT distance="675" swimtime="00:06:31.11" />
                    <SPLIT distance="700" swimtime="00:06:46.09" />
                    <SPLIT distance="725" swimtime="00:07:01.25" />
                    <SPLIT distance="750" swimtime="00:07:16.61" />
                    <SPLIT distance="775" swimtime="00:07:31.91" />
                    <SPLIT distance="800" swimtime="00:07:46.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124399" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="118566" reactiontime="+47" />
                    <RELAYPOSITION number="3" athleteid="129690" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="124394" reactiontime="+52" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Canada">
              <RESULTS>
                <RESULT eventid="134" place="4" lane="7" heat="1" swimtime="00:01:43.56" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.72" />
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                    <SPLIT distance="75" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:00:55.53" />
                    <SPLIT distance="125" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:19.93" />
                    <SPLIT distance="175" swimtime="00:01:31.11" />
                    <SPLIT distance="200" swimtime="00:01:43.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129652" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="118566" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="124174" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="124058" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="6" lane="5" heat="1" swimtime="00:01:46.16" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:26.10" />
                    <SPLIT distance="75" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:00:56.18" />
                    <SPLIT distance="125" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:21.70" />
                    <SPLIT distance="175" swimtime="00:01:33.42" />
                    <SPLIT distance="200" swimtime="00:01:46.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156529" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="118565" reactiontime="+37" />
                    <RELAYPOSITION number="3" athleteid="101207" reactiontime="+46" />
                    <RELAYPOSITION number="4" athleteid="124394" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Canada">
              <RESULTS>
                <RESULT eventid="111" place="3" lane="8" heat="1" swimtime="00:01:36.93" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.78" />
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                    <SPLIT distance="75" swimtime="00:00:37.15" />
                    <SPLIT distance="100" swimtime="00:00:51.66" />
                    <SPLIT distance="125" swimtime="00:01:01.50" />
                    <SPLIT distance="150" swimtime="00:01:13.78" />
                    <SPLIT distance="175" swimtime="00:01:24.85" />
                    <SPLIT distance="200" swimtime="00:01:36.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129652" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="124292" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="214502" reactiontime="+93" />
                    <RELAYPOSITION number="4" athleteid="124174" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="8" lane="7" heat="4" swimtime="00:01:39.01" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                    <SPLIT distance="75" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:00:51.99" />
                    <SPLIT distance="125" swimtime="00:01:02.09" />
                    <SPLIT distance="150" swimtime="00:01:14.40" />
                    <SPLIT distance="175" swimtime="00:01:26.21" />
                    <SPLIT distance="200" swimtime="00:01:39.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156529" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="124292" reactiontime="+26" />
                    <RELAYPOSITION number="3" athleteid="214502" reactiontime="+12" />
                    <RELAYPOSITION number="4" athleteid="124394" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Canada">
              <RESULTS>
                <RESULT eventid="35" place="-1" lane="5" heat="3" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Cayman Islands" shortname="CAY" code="CAY" nation="CAY" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154726" lastname="CROOKS" firstname="Jordan" gender="M" birthdate="2002-05-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.79" eventid="14" heat="6" lane="6">
                  <MEETINFO date="2022-06-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.20" eventid="31" heat="6" lane="3">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="6" lane="4" heat="1" heatid="10114" swimtime="00:00:45.77" reactiontime="+61" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.12" />
                    <SPLIT distance="50" swimtime="00:00:21.32" />
                    <SPLIT distance="75" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:00:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="1" lane="6" heat="6" heatid="60014" swimtime="00:00:45.61" reactiontime="+62" points="950">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:21.70" />
                    <SPLIT distance="75" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="1" lane="4" heat="2" heatid="20214" swimtime="00:00:45.55" reactiontime="+60" points="953">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:21.63" />
                    <SPLIT distance="75" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="131" place="1" lane="4" heat="1" heatid="10131" swimtime="00:00:20.46" reactiontime="+60" points="956">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.81" />
                    <SPLIT distance="50" swimtime="00:00:20.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="1" lane="3" heat="6" heatid="60031" swimtime="00:00:20.36" reactiontime="+59" points="970">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.80" />
                    <SPLIT distance="50" swimtime="00:00:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="1" lane="4" heat="2" heatid="20231" swimtime="00:00:20.31" reactiontime="+59" points="978">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.83" />
                    <SPLIT distance="50" swimtime="00:00:20.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195801" lastname="CROOKS" firstname="Jillian Janis Geohagan" gender="F" birthdate="2006-06-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.34" eventid="13" heat="5" lane="5">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.44" eventid="4" heat="3" lane="6">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="26" lane="5" heat="5" heatid="50013" swimtime="00:00:54.20" reactiontime="+63" points="796">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.92" />
                    <SPLIT distance="75" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:00:54.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="24" lane="6" heat="3" heatid="30004" swimtime="00:00:26.40" reactiontime="+60" points="787">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Congo" shortname="CGO" code="CGO" nation="CGO" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197094" lastname="DOUMA" firstname="Yann Emmanuel" gender="M" birthdate="1992-08-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="41" heat="1" lane="3" />
                <ENTRY entrytime="00:00:26.73" eventid="31" heat="3" lane="2">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="-1" lane="3" heat="1" heatid="10041" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="68" lane="2" heat="3" heatid="30031" swimtime="00:00:26.33" reactiontime="+77" points="448">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197008" lastname="BOBIMBO" firstname="Vanessa" gender="F" birthdate="1999-12-08">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="30" place="-1" lane="3" heat="1" heatid="10030" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Chile" shortname="CHI" code="CHI" nation="CHI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="130436" lastname="MARIN" firstname="Ines" gender="F" birthdate="2001-04-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.99" eventid="13" heat="5" lane="7">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:00.02" eventid="43" heat="2" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="35" lane="7" heat="5" heatid="50013" swimtime="00:00:55.28" reactiontime="+63" points="751">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                    <SPLIT distance="75" swimtime="00:00:40.88" />
                    <SPLIT distance="100" swimtime="00:00:55.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="22" lane="6" heat="2" heatid="20043" swimtime="00:01:58.79" reactiontime="+64" points="800">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="75" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:00:57.67" />
                    <SPLIT distance="125" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:27.93" />
                    <SPLIT distance="175" swimtime="00:01:43.58" />
                    <SPLIT distance="200" swimtime="00:01:58.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="China" shortname="CHN" code="CHN" nation="CHN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197625" lastname="WANG" firstname="Gukailai" gender="M" birthdate="2003-08-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.94" eventid="3" heat="5" lane="8">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.65" eventid="19" heat="5" lane="1">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="23" lane="8" heat="5" heatid="50003" swimtime="00:00:51.85" reactiontime="+58" points="809">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:24.89" />
                    <SPLIT distance="75" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:00:51.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="26" lane="1" heat="5" heatid="50019" swimtime="00:00:23.97" reactiontime="+55" points="796">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.81" />
                    <SPLIT distance="50" swimtime="00:00:23.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145336" lastname="QIN" firstname="Haiyang" gender="M" birthdate="1999-05-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.31" eventid="16" heat="7" lane="5">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.08" eventid="29" heat="4" lane="5">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.51" eventid="7" heat="5" lane="7">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:26.12" eventid="41" heat="7" lane="3">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="4" lane="3" heat="1" heatid="10116" swimtime="00:00:56.33" reactiontime="+63" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                    <SPLIT distance="75" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:00:56.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="3" lane="5" heat="7" heatid="70016" swimtime="00:00:56.66" reactiontime="+66" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.08" />
                    <SPLIT distance="50" swimtime="00:00:26.50" />
                    <SPLIT distance="75" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:00:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="3" lane="5" heat="2" heatid="20216" swimtime="00:00:56.38" reactiontime="+65" points="942">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="75" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:00:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="129" place="3" lane="6" heat="1" heatid="10129" swimtime="00:02:02.22" reactiontime="+66" points="950">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                    <SPLIT distance="125" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:01:30.22" />
                    <SPLIT distance="175" swimtime="00:01:46.26" />
                    <SPLIT distance="200" swimtime="00:02:02.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="4" lane="5" heat="4" heatid="40029" swimtime="00:02:03.81" reactiontime="+67" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="75" swimtime="00:00:43.22" />
                    <SPLIT distance="100" swimtime="00:00:59.14" />
                    <SPLIT distance="125" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:31.14" />
                    <SPLIT distance="175" swimtime="00:01:47.70" />
                    <SPLIT distance="200" swimtime="00:02:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="18" lane="7" heat="5" heatid="50007" swimtime="00:01:54.98" reactiontime="+66" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.96" />
                    <SPLIT distance="50" swimtime="00:00:24.48" />
                    <SPLIT distance="75" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:00:53.62" />
                    <SPLIT distance="125" swimtime="00:01:10.06" />
                    <SPLIT distance="150" swimtime="00:01:26.33" />
                    <SPLIT distance="175" swimtime="00:01:41.41" />
                    <SPLIT distance="200" swimtime="00:01:54.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="4" lane="7" heat="1" heatid="10141" swimtime="00:00:25.82" reactiontime="+65" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="5" lane="3" heat="7" heatid="70041" swimtime="00:00:26.13" reactiontime="+64" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="5" lane="3" heat="2" heatid="20241" swimtime="00:00:25.81" reactiontime="+63" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151731" lastname="SUN" firstname="Jiajun" gender="M" birthdate="2000-08-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.43" eventid="16" heat="6" lane="5">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.06" eventid="29" heat="5" lane="7">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="17" lane="5" heat="6" heatid="60016" swimtime="00:00:57.92" reactiontime="+69" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.37" />
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                    <SPLIT distance="75" swimtime="00:00:42.24" />
                    <SPLIT distance="100" swimtime="00:00:57.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="-1" lane="7" heat="5" heatid="50029" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201768" lastname="CHEN" firstname="Juner" gender="M" birthdate="2004-02-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.95" eventid="39" heat="8" lane="7">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:01:49.61" eventid="21" heat="2" lane="4">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:22.72" eventid="5" heat="8" lane="1">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="18" lane="7" heat="8" heatid="80039" swimtime="00:00:50.83" reactiontime="+64" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.77" />
                    <SPLIT distance="50" swimtime="00:00:23.54" />
                    <SPLIT distance="75" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:00:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="9" lane="4" heat="2" heatid="20021" swimtime="00:01:51.24" reactiontime="+62" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.32" />
                    <SPLIT distance="50" swimtime="00:00:25.59" />
                    <SPLIT distance="75" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:00:54.19" />
                    <SPLIT distance="125" swimtime="00:01:08.66" />
                    <SPLIT distance="150" swimtime="00:01:22.72" />
                    <SPLIT distance="175" swimtime="00:01:37.11" />
                    <SPLIT distance="200" swimtime="00:01:51.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="-1" lane="1" heat="8" heatid="80005" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197577" lastname="PAN" firstname="Zhanle" gender="M" birthdate="2004-08-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.27" eventid="14" heat="10" lane="5">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.66" eventid="44" heat="6" lane="2">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:53.10" eventid="23" heat="3" lane="7">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="6" lane="1" heat="1" heatid="10114" swimtime="00:00:45.77" reactiontime="+60" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.36" />
                    <SPLIT distance="50" swimtime="00:00:21.91" />
                    <SPLIT distance="75" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:00:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="11" lane="5" heat="10" heatid="100014" swimtime="00:00:46.79" reactiontime="+62" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.53" />
                    <SPLIT distance="75" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:00:46.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="7" lane="7" heat="2" heatid="20214" swimtime="00:00:46.19" reactiontime="+62" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.46" />
                    <SPLIT distance="50" swimtime="00:00:22.09" />
                    <SPLIT distance="75" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:00:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="14" lane="2" heat="6" heatid="60044" swimtime="00:01:43.48" reactiontime="+63" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.13" />
                    <SPLIT distance="50" swimtime="00:00:23.89" />
                    <SPLIT distance="75" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:00:50.49" />
                    <SPLIT distance="125" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:17.32" />
                    <SPLIT distance="175" swimtime="00:01:30.57" />
                    <SPLIT distance="200" swimtime="00:01:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="28" lane="7" heat="3" heatid="30023" swimtime="00:00:54.63" reactiontime="+63" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.07" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                    <SPLIT distance="75" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:00:54.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214429" lastname="WANG" firstname="Haoyu" gender="M" birthdate="2005-07-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.78" eventid="14" heat="11" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.77" eventid="31" heat="8" lane="1">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="24" lane="2" heat="11" heatid="110014" swimtime="00:00:47.17" reactiontime="+62" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.87" />
                    <SPLIT distance="50" swimtime="00:00:22.84" />
                    <SPLIT distance="75" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:00:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="37" lane="1" heat="8" heatid="80031" swimtime="00:00:21.60" reactiontime="+58" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:21.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191659" lastname="FEI" firstname="Liwei" gender="M" birthdate="2003-03-12">
              <ENTRIES>
                <ENTRY entrytime="00:14:35.50" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:03:41.56" eventid="24" heat="4" lane="8">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:07:37.74" eventid="42">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="-1" lane="7" heat="5" heatid="30110" swimtime="NT" status="DNS" />
                <RESULT eventid="24" place="-1" lane="8" heat="4" heatid="40024" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214430" lastname="TAO" firstname="Guannan" gender="M" birthdate="2004-04-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.75" eventid="46" heat="2" lane="7">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:04:17.13" eventid="37" heat="1" lane="6">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="15" lane="7" heat="2" heatid="20046" swimtime="00:01:53.14" reactiontime="+62" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="75" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:00:55.21" />
                    <SPLIT distance="125" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:24.04" />
                    <SPLIT distance="175" swimtime="00:01:38.67" />
                    <SPLIT distance="200" swimtime="00:01:53.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="19" lane="6" heat="1" heatid="10037" swimtime="00:04:14.85" reactiontime="+70" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.15" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:00:58.67" />
                    <SPLIT distance="125" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:30.92" />
                    <SPLIT distance="175" swimtime="00:01:47.17" />
                    <SPLIT distance="200" swimtime="00:02:02.87" />
                    <SPLIT distance="225" swimtime="00:02:21.02" />
                    <SPLIT distance="250" swimtime="00:02:39.58" />
                    <SPLIT distance="275" swimtime="00:02:57.48" />
                    <SPLIT distance="300" swimtime="00:03:15.89" />
                    <SPLIT distance="325" swimtime="00:03:31.87" />
                    <SPLIT distance="350" swimtime="00:03:46.94" />
                    <SPLIT distance="375" swimtime="00:04:01.49" />
                    <SPLIT distance="400" swimtime="00:04:14.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214428" lastname="XU" firstname="Fang" gender="M" birthdate="2003-05-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.52" eventid="21" heat="2" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="21" place="-1" lane="2" heat="2" heatid="20021" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214427" lastname="HUANG" firstname="Zhiwei" gender="M" birthdate="2000-07-10">
              <ENTRIES>
                <ENTRY entrytime="00:04:06.68" eventid="37" heat="2" lane="2">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="37" place="17" lane="2" heat="2" heatid="20037" swimtime="00:04:13.19" reactiontime="+68" points="797">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="75" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:00:55.63" />
                    <SPLIT distance="125" swimtime="00:01:11.64" />
                    <SPLIT distance="150" swimtime="00:01:27.28" />
                    <SPLIT distance="175" swimtime="00:01:42.94" />
                    <SPLIT distance="200" swimtime="00:01:58.50" />
                    <SPLIT distance="225" swimtime="00:02:16.48" />
                    <SPLIT distance="250" swimtime="00:02:35.04" />
                    <SPLIT distance="275" swimtime="00:02:53.75" />
                    <SPLIT distance="300" swimtime="00:03:12.83" />
                    <SPLIT distance="325" swimtime="00:03:28.55" />
                    <SPLIT distance="350" swimtime="00:03:43.48" />
                    <SPLIT distance="375" swimtime="00:03:58.80" />
                    <SPLIT distance="400" swimtime="00:04:13.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129462" lastname="YAN" firstname="Zibei" gender="M" birthdate="1995-10-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.16" eventid="41" heat="7" lane="6">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="141" place="7" lane="6" heat="1" heatid="10141" swimtime="00:00:26.06" reactiontime="+63" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="3" lane="6" heat="7" heatid="70041" swimtime="00:00:26.06" reactiontime="+61" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                    <SPLIT distance="50" swimtime="00:00:26.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="4" lane="5" heat="2" heatid="20241" swimtime="00:00:25.80" reactiontime="+61" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151732" lastname="PENG" firstname="Xuwei" gender="F" birthdate="2003-01-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.01" eventid="2" heat="4" lane="6">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.00" eventid="45" heat="4" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:26.56" eventid="18" heat="5" lane="7">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="17" lane="6" heat="4" heatid="40002" swimtime="00:00:57.67" reactiontime="+57" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="75" swimtime="00:00:42.83" />
                    <SPLIT distance="100" swimtime="00:00:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="6" lane="7" heat="1" heatid="10145" swimtime="00:02:02.39" reactiontime="+58" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                    <SPLIT distance="75" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:00:59.57" />
                    <SPLIT distance="125" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:31.14" />
                    <SPLIT distance="175" swimtime="00:01:46.95" />
                    <SPLIT distance="200" swimtime="00:02:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="6" lane="3" heat="4" heatid="40045" swimtime="00:02:03.27" reactiontime="+60" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="75" swimtime="00:00:44.24" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="125" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:31.78" />
                    <SPLIT distance="175" swimtime="00:01:47.75" />
                    <SPLIT distance="200" swimtime="00:02:03.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="22" lane="7" heat="5" heatid="50018" swimtime="00:00:26.99" reactiontime="+59" points="820">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:26.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197538" lastname="WAN" firstname="Letian" gender="F" birthdate="2004-08-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.05" eventid="2" heat="6" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:26.12" eventid="18" heat="6" lane="3">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="13" lane="2" heat="6" heatid="60002" swimtime="00:00:57.49" reactiontime="+56" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:42.42" />
                    <SPLIT distance="100" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="14" lane="1" heat="2" heatid="20202" swimtime="00:00:57.59" reactiontime="+57" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                    <SPLIT distance="75" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="12" lane="3" heat="6" heatid="60018" swimtime="00:00:26.38" reactiontime="+56" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="14" lane="7" heat="1" heatid="10218" swimtime="00:00:26.48" reactiontime="+55" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124144" lastname="YANG" firstname="Chang" gender="F" birthdate="2001-09-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.18" eventid="15" heat="7" lane="7">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.98" eventid="28" heat="3" lane="6">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="15" lane="7" heat="7" heatid="70015" swimtime="00:01:05.28" reactiontime="+68" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.16" />
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="75" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="11" lane="8" heat="1" heatid="10215" swimtime="00:01:04.99" reactiontime="+66" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="75" swimtime="00:00:47.48" />
                    <SPLIT distance="100" swimtime="00:01:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="22" lane="6" heat="3" heatid="30028" swimtime="00:02:24.80" reactiontime="+66" points="802">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.99" />
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="75" swimtime="00:00:50.80" />
                    <SPLIT distance="100" swimtime="00:01:08.77" />
                    <SPLIT distance="125" swimtime="00:01:27.24" />
                    <SPLIT distance="150" swimtime="00:01:45.91" />
                    <SPLIT distance="175" swimtime="00:02:05.32" />
                    <SPLIT distance="200" swimtime="00:02:24.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191700" lastname="TANG" firstname="Qianting" gender="F" birthdate="2004-03-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.15" eventid="15" heat="6" lane="4">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.65" eventid="28" heat="4" lane="5">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:29.19" eventid="40" heat="5" lane="4">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="4" lane="7" heat="1" heatid="10115" swimtime="00:01:04.06" reactiontime="+70" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.49" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:46.85" />
                    <SPLIT distance="100" swimtime="00:01:04.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="4" lane="4" heat="6" heatid="60015" swimtime="00:01:04.07" reactiontime="+72" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="75" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="5" lane="5" heat="1" heatid="10215" swimtime="00:01:04.36" reactiontime="+69" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="75" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="128" place="5" lane="2" heat="1" heatid="10128" swimtime="00:02:19.28" reactiontime="+69" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="75" swimtime="00:00:48.99" />
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                    <SPLIT distance="125" swimtime="00:01:24.83" />
                    <SPLIT distance="150" swimtime="00:01:43.17" />
                    <SPLIT distance="175" swimtime="00:02:01.23" />
                    <SPLIT distance="200" swimtime="00:02:19.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="4" lane="5" heat="4" heatid="40028" swimtime="00:02:19.57" reactiontime="+70" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.10" />
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="75" swimtime="00:00:49.13" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="125" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:01:42.92" />
                    <SPLIT distance="175" swimtime="00:02:01.15" />
                    <SPLIT distance="200" swimtime="00:02:19.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="4" lane="6" heat="1" heatid="10140" swimtime="00:00:29.22" reactiontime="+68" points="933">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="2" lane="4" heat="5" heatid="50040" swimtime="00:00:29.38" reactiontime="+66" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="4" lane="4" heat="1" heatid="10240" swimtime="00:00:29.28" reactiontime="+69" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110581" lastname="ZHANG" firstname="Yufei" gender="F" birthdate="1998-04-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.46" eventid="38" heat="4" lane="5">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:24.91" eventid="4" heat="6" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.82" eventid="30" heat="8" lane="5">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="-1" lane="5" heat="4" heatid="40038" swimtime="NT" status="DNS" />
                <RESULT eventid="104" place="3" lane="5" heat="1" heatid="10104" swimtime="00:00:24.71" reactiontime="+61" points="960">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.34" />
                    <SPLIT distance="50" swimtime="00:00:24.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="1" lane="5" heat="6" heatid="60004" swimtime="00:00:24.75" reactiontime="+63" points="955">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.33" />
                    <SPLIT distance="50" swimtime="00:00:24.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="2" lane="4" heat="2" heatid="20204" swimtime="00:00:24.79" reactiontime="+61" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.29" />
                    <SPLIT distance="50" swimtime="00:00:24.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="-1" lane="5" heat="8" heatid="80030" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152002" lastname="WANG" firstname="Yichun" gender="F" birthdate="2005-04-04">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:56.57" eventid="38" heat="4" lane="3">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.40" eventid="4" heat="6" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="-1" lane="3" heat="4" heatid="40038" swimtime="NT" status="DNS" />
                <RESULT eventid="4" place="6" lane="2" heat="6" heatid="60004" swimtime="00:00:25.28" reactiontime="+65" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.57" />
                    <SPLIT distance="50" swimtime="00:00:25.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="9" lane="3" heat="1" heatid="10204" swimtime="00:00:25.14" reactiontime="+68" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.57" />
                    <SPLIT distance="50" swimtime="00:00:25.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145348" lastname="WU" firstname="Qingfeng" gender="F" birthdate="2003-01-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.23" eventid="13" heat="7" lane="7">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:00:23.86" eventid="30" heat="8" lane="3">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="-1" lane="7" heat="7" heatid="70013" swimtime="NT" status="DNS" />
                <RESULT eventid="30" place="12" lane="3" heat="8" heatid="80030" swimtime="00:00:24.33" reactiontime="+67" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="11" lane="1" heat="2" heatid="20230" swimtime="00:00:24.21" reactiontime="+67" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197535" lastname="CHENG" firstname="Yujie" gender="F" birthdate="2005-09-22">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.57" eventid="13" heat="7" lane="6">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="13" lane="6" heat="7" heatid="70013" swimtime="00:00:53.03" reactiontime="+68" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:25.67" />
                    <SPLIT distance="75" swimtime="00:00:39.43" />
                    <SPLIT distance="100" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="14" lane="1" heat="2" heatid="20213" swimtime="00:00:52.90" reactiontime="+66" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:25.28" />
                    <SPLIT distance="75" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:00:52.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122811" lastname="LIU" firstname="Yaxin" gender="F" birthdate="1999-06-16">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.46" eventid="45" heat="4" lane="6">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:04:00.33" eventid="1" heat="3" lane="5">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="14" lane="6" heat="4" heatid="40045" swimtime="00:02:05.10" reactiontime="+63" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="75" swimtime="00:00:45.83" />
                    <SPLIT distance="100" swimtime="00:01:01.71" />
                    <SPLIT distance="125" swimtime="00:01:17.73" />
                    <SPLIT distance="150" swimtime="00:01:33.83" />
                    <SPLIT distance="175" swimtime="00:01:49.90" />
                    <SPLIT distance="200" swimtime="00:02:05.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="9" lane="5" heat="3" heatid="30001" swimtime="00:04:02.36" reactiontime="+75" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="75" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:00:58.59" />
                    <SPLIT distance="125" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:29.37" />
                    <SPLIT distance="175" swimtime="00:01:44.84" />
                    <SPLIT distance="200" swimtime="00:02:00.34" />
                    <SPLIT distance="225" swimtime="00:02:15.70" />
                    <SPLIT distance="250" swimtime="00:02:30.99" />
                    <SPLIT distance="275" swimtime="00:02:46.38" />
                    <SPLIT distance="300" swimtime="00:03:01.71" />
                    <SPLIT distance="325" swimtime="00:03:17.04" />
                    <SPLIT distance="350" swimtime="00:03:32.46" />
                    <SPLIT distance="375" swimtime="00:03:47.84" />
                    <SPLIT distance="400" swimtime="00:04:02.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214432" lastname="ZHANG" firstname="Yifan" gender="F" birthdate="2000-11-22">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.35" eventid="20" heat="4" lane="4">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="12" lane="4" heat="4" heatid="40020" swimtime="00:02:07.05" reactiontime="+68" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                    <SPLIT distance="75" swimtime="00:00:44.33" />
                    <SPLIT distance="100" swimtime="00:01:00.30" />
                    <SPLIT distance="125" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:01:33.10" />
                    <SPLIT distance="175" swimtime="00:01:50.19" />
                    <SPLIT distance="200" swimtime="00:02:07.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129468" lastname="LI" firstname="Bingjie" gender="F" birthdate="2002-03-03">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.25" eventid="43" heat="4" lane="4">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:03:51.30" eventid="1" heat="4" lane="4">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:15:41.80" eventid="33">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="-1" lane="4" heat="4" heatid="40043" swimtime="NT" status="DNS" />
                <RESULT eventid="1" place="-1" lane="4" heat="4" heatid="40001" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201767" lastname="GE" firstname="Chutong" gender="F" birthdate="2003-09-23">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.98" eventid="6" heat="2" lane="3">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="00:04:31.10" eventid="36" heat="3" lane="6">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="-1" lane="3" heat="2" heatid="20006" swimtime="NT" status="DNS" />
                <RESULT eventid="36" place="21" lane="6" heat="3" heatid="30036" swimtime="00:04:46.59" reactiontime="+74" points="737">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="75" swimtime="00:00:46.98" />
                    <SPLIT distance="100" swimtime="00:01:04.87" />
                    <SPLIT distance="125" swimtime="00:01:24.44" />
                    <SPLIT distance="150" swimtime="00:01:42.86" />
                    <SPLIT distance="175" swimtime="00:02:00.77" />
                    <SPLIT distance="200" swimtime="00:02:18.40" />
                    <SPLIT distance="225" swimtime="00:02:38.55" />
                    <SPLIT distance="250" swimtime="00:02:59.51" />
                    <SPLIT distance="275" swimtime="00:03:20.55" />
                    <SPLIT distance="300" swimtime="00:03:41.27" />
                    <SPLIT distance="325" swimtime="00:03:58.66" />
                    <SPLIT distance="350" swimtime="00:04:14.91" />
                    <SPLIT distance="375" swimtime="00:04:31.27" />
                    <SPLIT distance="400" swimtime="00:04:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165399" lastname="ZHANG" firstname="Ke" gender="F" birthdate="2001-04-12">
              <ENTRIES>
                <ENTRY entrytime="00:08:13.92" eventid="12" heat="0" lane="2147483647">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:15:52.30" eventid="33" heat="0" lane="2147483647">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="7" lane="3" heat="5" heatid="30112" swimtime="00:08:24.24" reactiontime="+66" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="75" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:00:59.59" />
                    <SPLIT distance="125" swimtime="00:01:15.03" />
                    <SPLIT distance="150" swimtime="00:01:30.57" />
                    <SPLIT distance="175" swimtime="00:01:46.11" />
                    <SPLIT distance="200" swimtime="00:02:01.60" />
                    <SPLIT distance="225" swimtime="00:02:17.06" />
                    <SPLIT distance="250" swimtime="00:02:32.57" />
                    <SPLIT distance="275" swimtime="00:02:48.16" />
                    <SPLIT distance="300" swimtime="00:03:03.72" />
                    <SPLIT distance="325" swimtime="00:03:19.38" />
                    <SPLIT distance="350" swimtime="00:03:34.98" />
                    <SPLIT distance="375" swimtime="00:03:50.74" />
                    <SPLIT distance="400" swimtime="00:04:06.40" />
                    <SPLIT distance="425" swimtime="00:04:22.11" />
                    <SPLIT distance="450" swimtime="00:04:37.83" />
                    <SPLIT distance="475" swimtime="00:04:53.56" />
                    <SPLIT distance="500" swimtime="00:05:09.27" />
                    <SPLIT distance="525" swimtime="00:05:25.05" />
                    <SPLIT distance="550" swimtime="00:05:40.79" />
                    <SPLIT distance="575" swimtime="00:05:56.78" />
                    <SPLIT distance="600" swimtime="00:06:12.62" />
                    <SPLIT distance="625" swimtime="00:06:28.62" />
                    <SPLIT distance="650" swimtime="00:06:44.72" />
                    <SPLIT distance="675" swimtime="00:07:01.22" />
                    <SPLIT distance="700" swimtime="00:07:17.73" />
                    <SPLIT distance="725" swimtime="00:07:34.51" />
                    <SPLIT distance="750" swimtime="00:07:51.08" />
                    <SPLIT distance="775" swimtime="00:08:08.09" />
                    <SPLIT distance="800" swimtime="00:08:24.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="4" lane="6" heat="5" heatid="30133" swimtime="00:15:51.64" reactiontime="+66" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="75" swimtime="00:00:44.82" />
                    <SPLIT distance="100" swimtime="00:01:00.76" />
                    <SPLIT distance="125" swimtime="00:01:16.70" />
                    <SPLIT distance="150" swimtime="00:01:32.68" />
                    <SPLIT distance="175" swimtime="00:01:48.50" />
                    <SPLIT distance="200" swimtime="00:02:04.54" />
                    <SPLIT distance="225" swimtime="00:02:20.31" />
                    <SPLIT distance="250" swimtime="00:02:36.20" />
                    <SPLIT distance="275" swimtime="00:02:52.12" />
                    <SPLIT distance="300" swimtime="00:03:08.29" />
                    <SPLIT distance="325" swimtime="00:03:24.25" />
                    <SPLIT distance="350" swimtime="00:03:40.20" />
                    <SPLIT distance="375" swimtime="00:03:56.10" />
                    <SPLIT distance="400" swimtime="00:04:11.94" />
                    <SPLIT distance="425" swimtime="00:04:27.86" />
                    <SPLIT distance="450" swimtime="00:04:43.84" />
                    <SPLIT distance="475" swimtime="00:04:59.85" />
                    <SPLIT distance="500" swimtime="00:05:15.68" />
                    <SPLIT distance="525" swimtime="00:05:31.70" />
                    <SPLIT distance="550" swimtime="00:05:47.56" />
                    <SPLIT distance="575" swimtime="00:06:03.64" />
                    <SPLIT distance="600" swimtime="00:06:19.52" />
                    <SPLIT distance="625" swimtime="00:06:35.59" />
                    <SPLIT distance="650" swimtime="00:06:51.52" />
                    <SPLIT distance="675" swimtime="00:07:07.61" />
                    <SPLIT distance="700" swimtime="00:07:23.57" />
                    <SPLIT distance="725" swimtime="00:07:39.74" />
                    <SPLIT distance="750" swimtime="00:07:55.90" />
                    <SPLIT distance="775" swimtime="00:08:11.83" />
                    <SPLIT distance="800" swimtime="00:08:27.77" />
                    <SPLIT distance="825" swimtime="00:08:43.75" />
                    <SPLIT distance="850" swimtime="00:08:59.65" />
                    <SPLIT distance="875" swimtime="00:09:15.73" />
                    <SPLIT distance="900" swimtime="00:09:31.68" />
                    <SPLIT distance="925" swimtime="00:09:47.74" />
                    <SPLIT distance="950" swimtime="00:10:03.79" />
                    <SPLIT distance="975" swimtime="00:10:19.93" />
                    <SPLIT distance="1000" swimtime="00:10:35.78" />
                    <SPLIT distance="1025" swimtime="00:10:51.89" />
                    <SPLIT distance="1050" swimtime="00:11:07.86" />
                    <SPLIT distance="1075" swimtime="00:11:23.92" />
                    <SPLIT distance="1100" swimtime="00:11:39.73" />
                    <SPLIT distance="1125" swimtime="00:11:55.76" />
                    <SPLIT distance="1150" swimtime="00:12:11.65" />
                    <SPLIT distance="1175" swimtime="00:12:27.73" />
                    <SPLIT distance="1200" swimtime="00:12:43.53" />
                    <SPLIT distance="1225" swimtime="00:12:59.58" />
                    <SPLIT distance="1250" swimtime="00:13:15.44" />
                    <SPLIT distance="1275" swimtime="00:13:31.39" />
                    <SPLIT distance="1300" swimtime="00:13:47.16" />
                    <SPLIT distance="1325" swimtime="00:14:03.17" />
                    <SPLIT distance="1350" swimtime="00:14:18.92" />
                    <SPLIT distance="1375" swimtime="00:14:34.89" />
                    <SPLIT distance="1400" swimtime="00:14:50.64" />
                    <SPLIT distance="1425" swimtime="00:15:06.45" />
                    <SPLIT distance="1450" swimtime="00:15:22.15" />
                    <SPLIT distance="1475" swimtime="00:15:37.32" />
                    <SPLIT distance="1500" swimtime="00:15:51.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197578" lastname="CHEN" firstname="Ende" gender="M" birthdate="2004-04-07" />
            <ATHLETE athleteid="214431" lastname="LIU" firstname="Shuhan" gender="F" birthdate="2006-01-29" />
            <ATHLETE athleteid="145364" lastname="YANG" firstname="Junxuan" gender="F" birthdate="2002-01-26" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="9" place="-1" lane="3" heat="2" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="148" place="7" lane="1" heat="1" swimtime="00:03:25.15" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:24.56" />
                    <SPLIT distance="75" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:00:51.54" />
                    <SPLIT distance="125" swimtime="00:01:03.62" />
                    <SPLIT distance="150" swimtime="00:01:17.96" />
                    <SPLIT distance="175" swimtime="00:01:33.15" />
                    <SPLIT distance="200" swimtime="00:01:48.90" />
                    <SPLIT distance="225" swimtime="00:01:59.07" />
                    <SPLIT distance="250" swimtime="00:02:11.44" />
                    <SPLIT distance="275" swimtime="00:02:25.05" />
                    <SPLIT distance="300" swimtime="00:02:39.06" />
                    <SPLIT distance="325" swimtime="00:02:49.24" />
                    <SPLIT distance="350" swimtime="00:03:01.18" />
                    <SPLIT distance="375" swimtime="00:03:13.12" />
                    <SPLIT distance="400" swimtime="00:03:25.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197625" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="145336" reactiontime="+49" />
                    <RELAYPOSITION number="3" athleteid="201768" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="197577" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="7" lane="2" heat="2" swimtime="00:03:26.01" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:25.05" />
                    <SPLIT distance="75" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:00:51.82" />
                    <SPLIT distance="125" swimtime="00:01:04.04" />
                    <SPLIT distance="150" swimtime="00:01:18.80" />
                    <SPLIT distance="175" swimtime="00:01:33.95" />
                    <SPLIT distance="200" swimtime="00:01:49.43" />
                    <SPLIT distance="225" swimtime="00:01:59.94" />
                    <SPLIT distance="250" swimtime="00:02:12.79" />
                    <SPLIT distance="275" swimtime="00:02:26.08" />
                    <SPLIT distance="300" swimtime="00:02:39.73" />
                    <SPLIT distance="325" swimtime="00:02:49.96" />
                    <SPLIT distance="350" swimtime="00:03:01.77" />
                    <SPLIT distance="375" swimtime="00:03:13.88" />
                    <SPLIT distance="400" swimtime="00:03:26.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197625" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="145336" reactiontime="+54" />
                    <RELAYPOSITION number="3" athleteid="201768" reactiontime="+42" />
                    <RELAYPOSITION number="4" athleteid="197577" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="32" place="11" lane="5" heat="1" swimtime="00:07:06.26" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:24.31" />
                    <SPLIT distance="75" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:00:51.48" />
                    <SPLIT distance="125" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:18.24" />
                    <SPLIT distance="175" swimtime="00:01:31.87" />
                    <SPLIT distance="200" swimtime="00:01:44.85" />
                    <SPLIT distance="225" swimtime="00:01:55.77" />
                    <SPLIT distance="250" swimtime="00:02:08.56" />
                    <SPLIT distance="275" swimtime="00:02:21.94" />
                    <SPLIT distance="300" swimtime="00:02:35.59" />
                    <SPLIT distance="325" swimtime="00:02:49.53" />
                    <SPLIT distance="350" swimtime="00:03:03.51" />
                    <SPLIT distance="375" swimtime="00:03:17.41" />
                    <SPLIT distance="400" swimtime="00:03:30.89" />
                    <SPLIT distance="425" swimtime="00:03:41.83" />
                    <SPLIT distance="450" swimtime="00:03:54.80" />
                    <SPLIT distance="475" swimtime="00:04:08.15" />
                    <SPLIT distance="500" swimtime="00:04:21.76" />
                    <SPLIT distance="525" swimtime="00:04:35.22" />
                    <SPLIT distance="550" swimtime="00:04:48.94" />
                    <SPLIT distance="575" swimtime="00:05:02.78" />
                    <SPLIT distance="600" swimtime="00:05:16.22" />
                    <SPLIT distance="625" swimtime="00:05:27.58" />
                    <SPLIT distance="650" swimtime="00:05:40.42" />
                    <SPLIT distance="675" swimtime="00:05:54.17" />
                    <SPLIT distance="700" swimtime="00:06:08.08" />
                    <SPLIT distance="725" swimtime="00:06:22.26" />
                    <SPLIT distance="750" swimtime="00:06:36.93" />
                    <SPLIT distance="775" swimtime="00:06:51.73" />
                    <SPLIT distance="800" swimtime="00:07:06.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197577" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="214430" reactiontime="+14" />
                    <RELAYPOSITION number="3" athleteid="201768" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="197578" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="26" place="-1" lane="5" heat="1" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="127" place="6" lane="2" heat="1" swimtime="00:01:30.18" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.40" />
                    <SPLIT distance="50" swimtime="00:00:21.49" />
                    <SPLIT distance="75" swimtime="00:00:31.30" />
                    <SPLIT distance="100" swimtime="00:00:42.38" />
                    <SPLIT distance="125" swimtime="00:00:53.60" />
                    <SPLIT distance="150" swimtime="00:01:06.36" />
                    <SPLIT distance="175" swimtime="00:01:17.55" />
                    <SPLIT distance="200" swimtime="00:01:30.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197577" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="214429" reactiontime="+6" />
                    <RELAYPOSITION number="3" athleteid="152002" reactiontime="+10" />
                    <RELAYPOSITION number="4" athleteid="214431" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="5" lane="7" heat="3" swimtime="00:01:31.21" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.44" />
                    <SPLIT distance="50" swimtime="00:00:21.53" />
                    <SPLIT distance="75" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:00:42.67" />
                    <SPLIT distance="125" swimtime="00:00:54.34" />
                    <SPLIT distance="150" swimtime="00:01:07.03" />
                    <SPLIT distance="175" swimtime="00:01:18.60" />
                    <SPLIT distance="200" swimtime="00:01:31.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197577" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="214429" reactiontime="+6" />
                    <RELAYPOSITION number="3" athleteid="152002" reactiontime="+40" />
                    <RELAYPOSITION number="4" athleteid="214431" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="108" place="6" lane="2" heat="1" swimtime="00:03:29.96" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:25.37" />
                    <SPLIT distance="75" swimtime="00:00:39.24" />
                    <SPLIT distance="100" swimtime="00:00:53.02" />
                    <SPLIT distance="125" swimtime="00:01:04.65" />
                    <SPLIT distance="150" swimtime="00:01:18.02" />
                    <SPLIT distance="175" swimtime="00:01:31.92" />
                    <SPLIT distance="200" swimtime="00:01:45.53" />
                    <SPLIT distance="225" swimtime="00:01:57.21" />
                    <SPLIT distance="250" swimtime="00:02:10.61" />
                    <SPLIT distance="275" swimtime="00:02:24.37" />
                    <SPLIT distance="300" swimtime="00:02:38.05" />
                    <SPLIT distance="325" swimtime="00:02:49.08" />
                    <SPLIT distance="350" swimtime="00:03:02.45" />
                    <SPLIT distance="375" swimtime="00:03:16.51" />
                    <SPLIT distance="400" swimtime="00:03:29.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="145364" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="197535" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="145348" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="110581" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="5" lane="3" heat="1" swimtime="00:03:32.05" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.03" />
                    <SPLIT distance="50" swimtime="00:00:25.41" />
                    <SPLIT distance="75" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:00:52.95" />
                    <SPLIT distance="125" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:18.18" />
                    <SPLIT distance="175" swimtime="00:01:32.17" />
                    <SPLIT distance="200" swimtime="00:01:45.89" />
                    <SPLIT distance="225" swimtime="00:01:57.85" />
                    <SPLIT distance="250" swimtime="00:02:11.28" />
                    <SPLIT distance="275" swimtime="00:02:25.24" />
                    <SPLIT distance="300" swimtime="00:02:38.85" />
                    <SPLIT distance="325" swimtime="00:02:50.81" />
                    <SPLIT distance="350" swimtime="00:03:04.36" />
                    <SPLIT distance="375" swimtime="00:03:18.39" />
                    <SPLIT distance="400" swimtime="00:03:32.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="145364" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="214431" reactiontime="+35" />
                    <RELAYPOSITION number="3" athleteid="145348" reactiontime="+45" />
                    <RELAYPOSITION number="4" athleteid="197535" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="147" place="7" lane="8" heat="1" swimtime="00:03:51.44" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:00:57.64" />
                    <SPLIT distance="125" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:26.94" />
                    <SPLIT distance="175" swimtime="00:01:43.79" />
                    <SPLIT distance="200" swimtime="00:02:01.20" />
                    <SPLIT distance="225" swimtime="00:02:13.14" />
                    <SPLIT distance="250" swimtime="00:02:27.72" />
                    <SPLIT distance="275" swimtime="00:02:43.01" />
                    <SPLIT distance="300" swimtime="00:02:58.69" />
                    <SPLIT distance="325" swimtime="00:03:10.25" />
                    <SPLIT distance="350" swimtime="00:03:23.55" />
                    <SPLIT distance="375" swimtime="00:03:37.44" />
                    <SPLIT distance="400" swimtime="00:03:51.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="151732" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="191700" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="145364" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="214431" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="8" lane="5" heat="2" swimtime="00:03:54.57" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.21" />
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="75" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:00:58.08" />
                    <SPLIT distance="125" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:29.00" />
                    <SPLIT distance="175" swimtime="00:01:45.85" />
                    <SPLIT distance="200" swimtime="00:02:03.34" />
                    <SPLIT distance="225" swimtime="00:02:15.30" />
                    <SPLIT distance="250" swimtime="00:02:29.91" />
                    <SPLIT distance="275" swimtime="00:02:45.17" />
                    <SPLIT distance="300" swimtime="00:03:00.66" />
                    <SPLIT distance="325" swimtime="00:03:12.84" />
                    <SPLIT distance="350" swimtime="00:03:26.47" />
                    <SPLIT distance="375" swimtime="00:03:40.65" />
                    <SPLIT distance="400" swimtime="00:03:54.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197538" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="124144" reactiontime="+52" />
                    <RELAYPOSITION number="3" athleteid="145364" reactiontime="+16" />
                    <RELAYPOSITION number="4" athleteid="197535" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="117" place="6" lane="6" heat="1" swimtime="00:07:48.73" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="75" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:00:56.90" />
                    <SPLIT distance="125" swimtime="00:01:11.20" />
                    <SPLIT distance="150" swimtime="00:01:25.81" />
                    <SPLIT distance="175" swimtime="00:01:40.44" />
                    <SPLIT distance="200" swimtime="00:01:54.62" />
                    <SPLIT distance="225" swimtime="00:02:06.90" />
                    <SPLIT distance="250" swimtime="00:02:21.52" />
                    <SPLIT distance="275" swimtime="00:02:36.22" />
                    <SPLIT distance="300" swimtime="00:02:51.16" />
                    <SPLIT distance="325" swimtime="00:03:06.17" />
                    <SPLIT distance="350" swimtime="00:03:21.45" />
                    <SPLIT distance="375" swimtime="00:03:36.74" />
                    <SPLIT distance="400" swimtime="00:03:51.40" />
                    <SPLIT distance="425" swimtime="00:04:04.38" />
                    <SPLIT distance="450" swimtime="00:04:18.77" />
                    <SPLIT distance="475" swimtime="00:04:33.95" />
                    <SPLIT distance="500" swimtime="00:04:49.23" />
                    <SPLIT distance="525" swimtime="00:05:04.88" />
                    <SPLIT distance="550" swimtime="00:05:20.72" />
                    <SPLIT distance="575" swimtime="00:05:36.16" />
                    <SPLIT distance="600" swimtime="00:05:51.09" />
                    <SPLIT distance="625" swimtime="00:06:03.75" />
                    <SPLIT distance="650" swimtime="00:06:18.70" />
                    <SPLIT distance="675" swimtime="00:06:33.59" />
                    <SPLIT distance="700" swimtime="00:06:48.55" />
                    <SPLIT distance="725" swimtime="00:07:03.72" />
                    <SPLIT distance="750" swimtime="00:07:18.91" />
                    <SPLIT distance="775" swimtime="00:07:34.22" />
                    <SPLIT distance="800" swimtime="00:07:48.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="122811" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="145348" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="197535" reactiontime="+46" />
                    <RELAYPOSITION number="4" athleteid="214432" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="4" lane="5" heat="1" swimtime="00:07:45.88" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.50" />
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                    <SPLIT distance="75" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:00:56.12" />
                    <SPLIT distance="125" swimtime="00:01:11.09" />
                    <SPLIT distance="150" swimtime="00:01:26.72" />
                    <SPLIT distance="175" swimtime="00:01:42.54" />
                    <SPLIT distance="200" swimtime="00:01:57.89" />
                    <SPLIT distance="225" swimtime="00:02:10.37" />
                    <SPLIT distance="250" swimtime="00:02:24.81" />
                    <SPLIT distance="275" swimtime="00:02:39.94" />
                    <SPLIT distance="300" swimtime="00:02:55.31" />
                    <SPLIT distance="325" swimtime="00:03:10.41" />
                    <SPLIT distance="350" swimtime="00:03:25.69" />
                    <SPLIT distance="375" swimtime="00:03:41.22" />
                    <SPLIT distance="400" swimtime="00:03:55.88" />
                    <SPLIT distance="425" swimtime="00:04:08.29" />
                    <SPLIT distance="450" swimtime="00:04:22.56" />
                    <SPLIT distance="475" swimtime="00:04:37.25" />
                    <SPLIT distance="500" swimtime="00:04:51.74" />
                    <SPLIT distance="525" swimtime="00:05:06.09" />
                    <SPLIT distance="550" swimtime="00:05:20.54" />
                    <SPLIT distance="575" swimtime="00:05:35.42" />
                    <SPLIT distance="600" swimtime="00:05:49.78" />
                    <SPLIT distance="625" swimtime="00:06:02.37" />
                    <SPLIT distance="650" swimtime="00:06:16.96" />
                    <SPLIT distance="675" swimtime="00:06:31.58" />
                    <SPLIT distance="700" swimtime="00:06:46.27" />
                    <SPLIT distance="725" swimtime="00:07:01.18" />
                    <SPLIT distance="750" swimtime="00:07:16.24" />
                    <SPLIT distance="775" swimtime="00:07:31.40" />
                    <SPLIT distance="800" swimtime="00:07:45.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="145348" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="197535" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="122811" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="214432" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="125" place="5" lane="4" heat="1" swimtime="00:01:36.12" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:24.24" />
                    <SPLIT distance="75" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:00:47.91" />
                    <SPLIT distance="125" swimtime="00:00:59.34" />
                    <SPLIT distance="150" swimtime="00:01:11.97" />
                    <SPLIT distance="175" swimtime="00:01:23.49" />
                    <SPLIT distance="200" swimtime="00:01:36.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="145364" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="197535" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="214431" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="152002" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="1" lane="5" heat="1" swimtime="00:01:36.08" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:23.76" />
                    <SPLIT distance="75" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:00:47.82" />
                    <SPLIT distance="125" swimtime="00:00:59.47" />
                    <SPLIT distance="150" swimtime="00:01:11.92" />
                    <SPLIT distance="175" swimtime="00:01:23.61" />
                    <SPLIT distance="200" swimtime="00:01:36.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="110581" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="214431" reactiontime="+26" />
                    <RELAYPOSITION number="3" athleteid="197535" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="145364" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="34" place="10" lane="3" heat="2" swimtime="00:01:48.32" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                    <SPLIT distance="125" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:24.21" />
                    <SPLIT distance="175" swimtime="00:01:35.76" />
                    <SPLIT distance="200" swimtime="00:01:48.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="151732" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="124144" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="214432" reactiontime="+33" />
                    <RELAYPOSITION number="4" athleteid="214431" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="111" place="5" lane="1" heat="1" swimtime="00:01:37.31" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.67" />
                    <SPLIT distance="50" swimtime="00:00:23.74" />
                    <SPLIT distance="75" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:00:49.15" />
                    <SPLIT distance="125" swimtime="00:01:00.18" />
                    <SPLIT distance="150" swimtime="00:01:13.69" />
                    <SPLIT distance="175" swimtime="00:01:24.89" />
                    <SPLIT distance="200" swimtime="00:01:37.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197625" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="129462" reactiontime="+14" />
                    <RELAYPOSITION number="3" athleteid="110581" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="145348" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="7" lane="1" heat="1" swimtime="00:01:39.00" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                    <SPLIT distance="75" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:00:49.87" />
                    <SPLIT distance="125" swimtime="00:01:01.14" />
                    <SPLIT distance="150" swimtime="00:01:14.95" />
                    <SPLIT distance="175" swimtime="00:01:26.19" />
                    <SPLIT distance="200" swimtime="00:01:39.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197625" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="145336" reactiontime="+39" />
                    <RELAYPOSITION number="3" athleteid="152002" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="145348" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="People's Republic of China">
              <RESULTS>
                <RESULT eventid="135" place="7" lane="8" heat="1" swimtime="00:01:33.13" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:24.01" />
                    <SPLIT distance="75" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:00:49.73" />
                    <SPLIT distance="125" swimtime="00:00:59.90" />
                    <SPLIT distance="150" swimtime="00:01:12.25" />
                    <SPLIT distance="175" swimtime="00:01:22.15" />
                    <SPLIT distance="200" swimtime="00:01:33.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197625" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="129462" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="201768" reactiontime="+43" />
                    <RELAYPOSITION number="4" athleteid="197577" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="8" lane="3" heat="1" swimtime="00:01:34.24" reactiontime="+52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="75" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:00:50.06" />
                    <SPLIT distance="125" swimtime="00:01:00.16" />
                    <SPLIT distance="150" swimtime="00:01:12.58" />
                    <SPLIT distance="175" swimtime="00:01:23.00" />
                    <SPLIT distance="200" swimtime="00:01:34.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197625" reactiontime="+52" />
                    <RELAYPOSITION number="2" athleteid="145336" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="201768" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="214429" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Cameroon" shortname="CMR" code="CMR" nation="CMR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197184" lastname="NGUICHIE" firstname="Hugo Giovani" gender="M" birthdate="2007-07-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.63" eventid="14" heat="1" lane="3">
                  <MEETINFO date="2021-10-13" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.55" eventid="31" heat="2" lane="7">
                  <MEETINFO date="2021-10-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="-1" lane="3" heat="1" heatid="10014" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="-1" lane="7" heat="2" heatid="20031" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213128" lastname="ZENON" firstname="Cassandre  Athenais" gender="F" birthdate="2000-09-08">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="4" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="30" heat="2" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="34" lane="4" heat="1" heatid="10004" swimtime="00:00:29.32" reactiontime="+76" points="574">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="42" lane="1" heat="2" heatid="20030" swimtime="00:00:27.87" reactiontime="+73" points="556">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Cook Islands" shortname="COK" code="COK" nation="COK" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="128651" lastname="ROBERTS" firstname="Wesley Tikiariki" gender="M" birthdate="1997-06-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.39" eventid="14" heat="5" lane="5">
                  <MEETINFO date="2022-05-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.33" eventid="44" heat="2" lane="4">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:03:55.65" eventid="24" heat="2" lane="8">
                  <MEETINFO date="2021-07-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="47" lane="5" heat="5" heatid="50014" swimtime="00:00:49.59" reactiontime="+71" points="739">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.20" />
                    <SPLIT distance="50" swimtime="00:00:23.51" />
                    <SPLIT distance="75" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:00:49.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="29" lane="4" heat="2" heatid="20044" swimtime="00:01:46.67" reactiontime="+73" points="808">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:25.06" />
                    <SPLIT distance="75" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:00:52.23" />
                    <SPLIT distance="125" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:19.46" />
                    <SPLIT distance="175" swimtime="00:01:33.24" />
                    <SPLIT distance="200" swimtime="00:01:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="26" lane="8" heat="2" heatid="20024" swimtime="00:03:50.03" reactiontime="+74" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                    <SPLIT distance="75" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:00:54.18" />
                    <SPLIT distance="125" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:23.30" />
                    <SPLIT distance="175" swimtime="00:01:38.03" />
                    <SPLIT distance="200" swimtime="00:01:52.84" />
                    <SPLIT distance="225" swimtime="00:02:07.60" />
                    <SPLIT distance="250" swimtime="00:02:22.17" />
                    <SPLIT distance="275" swimtime="00:02:36.72" />
                    <SPLIT distance="300" swimtime="00:02:51.38" />
                    <SPLIT distance="325" swimtime="00:03:06.11" />
                    <SPLIT distance="350" swimtime="00:03:20.95" />
                    <SPLIT distance="375" swimtime="00:03:35.82" />
                    <SPLIT distance="400" swimtime="00:03:50.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140885" lastname="AITU" firstname="Bede" gender="M" birthdate="2001-10-11">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.49" eventid="46" heat="1" lane="2">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="-1" lane="2" heat="1" heatid="10046" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195483" lastname="CONNOLLY" firstname="Mary Lanihei" gender="F" birthdate="2005-12-30">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.76" eventid="15" heat="3" lane="1">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.77" eventid="40" heat="3" lane="4">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="34" lane="1" heat="3" heatid="30015" swimtime="00:01:07.66" reactiontime="+69" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.56" />
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="75" swimtime="00:00:49.49" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="27" lane="4" heat="3" heatid="30040" swimtime="00:00:31.68" reactiontime="+65" points="732">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.59" />
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129166" lastname="FISHER-MARSTERS" firstname="Kirsten Andrea" gender="F" birthdate="1998-02-11">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="6" heat="1" lane="3" />
                <ENTRY entrytime="00:01:06.67" eventid="22" heat="2" lane="8">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="34" lane="3" heat="1" heatid="10006" swimtime="00:02:28.89" reactiontime="+65" points="548">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="75" swimtime="00:00:50.39" />
                    <SPLIT distance="100" swimtime="00:01:09.08" />
                    <SPLIT distance="125" swimtime="00:01:30.11" />
                    <SPLIT distance="150" swimtime="00:01:51.43" />
                    <SPLIT distance="175" swimtime="00:02:11.22" />
                    <SPLIT distance="200" swimtime="00:02:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="26" lane="8" heat="2" heatid="20022" swimtime="00:01:07.40" reactiontime="+66" points="589">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.67" />
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="75" swimtime="00:00:50.03" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Colombia" shortname="COL" code="COL" nation="COL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="102352" lastname="MURILLO VALDES" firstname="Jorge" gender="M" birthdate="1991-09-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.58" eventid="16" heat="4" lane="1">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.46" eventid="29" heat="2" lane="1">
                  <MEETINFO date="2021-07-27" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.19" eventid="41" heat="6" lane="1">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="31" lane="1" heat="4" heatid="40016" swimtime="00:00:58.83" reactiontime="+63" points="829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                    <SPLIT distance="50" swimtime="00:00:27.59" />
                    <SPLIT distance="75" swimtime="00:00:42.96" />
                    <SPLIT distance="100" swimtime="00:00:58.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="23" lane="1" heat="2" heatid="20029" swimtime="00:02:08.91" reactiontime="+63" points="809">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="75" swimtime="00:00:44.72" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="125" swimtime="00:01:17.79" />
                    <SPLIT distance="150" swimtime="00:01:34.78" />
                    <SPLIT distance="175" swimtime="00:01:51.80" />
                    <SPLIT distance="200" swimtime="00:02:08.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="-1" lane="1" heat="6" heatid="60041" swimtime="00:00:27.09" status="DSQ" reactiontime="+65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125185" lastname="CORREDOR" firstname="Santiago" gender="M" birthdate="1999-05-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.80" eventid="44" heat="2" lane="2">
                  <MEETINFO date="2021-11-26" />
                </ENTRY>
                <ENTRY entrytime="00:03:47.53" eventid="24" heat="2" lane="5">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="32" lane="2" heat="2" heatid="20044" swimtime="00:01:47.47" reactiontime="+68" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:25.42" />
                    <SPLIT distance="75" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:00:52.61" />
                    <SPLIT distance="125" swimtime="00:01:05.99" />
                    <SPLIT distance="150" swimtime="00:01:19.70" />
                    <SPLIT distance="175" swimtime="00:01:33.79" />
                    <SPLIT distance="200" swimtime="00:01:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="22" lane="5" heat="2" heatid="20024" swimtime="00:03:47.60" reactiontime="+66" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:54.29" />
                    <SPLIT distance="125" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:22.52" />
                    <SPLIT distance="175" swimtime="00:01:36.88" />
                    <SPLIT distance="200" swimtime="00:01:51.19" />
                    <SPLIT distance="225" swimtime="00:02:05.66" />
                    <SPLIT distance="250" swimtime="00:02:20.17" />
                    <SPLIT distance="275" swimtime="00:02:34.82" />
                    <SPLIT distance="300" swimtime="00:02:49.25" />
                    <SPLIT distance="325" swimtime="00:03:03.68" />
                    <SPLIT distance="350" swimtime="00:03:18.29" />
                    <SPLIT distance="375" swimtime="00:03:33.15" />
                    <SPLIT distance="400" swimtime="00:03:47.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214514" lastname="GOMEZ HURTADO" firstname="Stefania" gender="F" birthdate="2004-04-12">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:08.49" eventid="15" heat="3" lane="4">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.63" eventid="22" heat="4" lane="7">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="35" lane="4" heat="3" heatid="30015" swimtime="00:01:08.71" reactiontime="+65" points="747">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.99" />
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="75" swimtime="00:00:50.18" />
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="18" lane="7" heat="4" heatid="40022" swimtime="00:01:01.27" reactiontime="+67" points="784">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                    <SPLIT distance="75" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:01.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156156" lastname="ROWE CERVANTES" firstname="Sirena Carolina" gender="F" birthdate="1998-02-28">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:26.42" eventid="4" heat="4" lane="1">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.00" eventid="30" heat="6" lane="8">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="22" lane="1" heat="4" heatid="40004" swimtime="00:00:26.12" reactiontime="+66" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="27" lane="8" heat="6" heatid="60030" swimtime="00:00:25.19" reactiontime="+68" points="754">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:25.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Colombia">
              <RESULTS>
                <RESULT eventid="27" place="14" lane="5" heat="1" swimtime="00:01:35.07" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.21" />
                    <SPLIT distance="50" swimtime="00:00:22.99" />
                    <SPLIT distance="75" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:00:45.77" />
                    <SPLIT distance="125" swimtime="00:00:57.55" />
                    <SPLIT distance="150" swimtime="00:01:10.83" />
                    <SPLIT distance="175" swimtime="00:01:22.21" />
                    <SPLIT distance="200" swimtime="00:01:35.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="125185" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="102352" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="214514" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="156156" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Colombia">
              <RESULTS>
                <RESULT eventid="11" place="16" lane="2" heat="2" swimtime="00:01:42.46" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:24.77" />
                    <SPLIT distance="75" swimtime="00:00:36.48" />
                    <SPLIT distance="100" swimtime="00:00:51.26" />
                    <SPLIT distance="125" swimtime="00:01:02.78" />
                    <SPLIT distance="150" swimtime="00:01:17.42" />
                    <SPLIT distance="175" swimtime="00:01:29.25" />
                    <SPLIT distance="200" swimtime="00:01:42.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="125185" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="102352" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="156156" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="214514" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Comoros" shortname="COM" code="COM" nation="COM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="164063" lastname="MOHAMED" firstname="Ibrahim" gender="M" birthdate="1996-01-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.58" eventid="5" heat="2" lane="4">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="-1" lane="4" heat="2" heatid="20005" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156558" lastname="YOUSSOUF" firstname="Hakim" gender="M" birthdate="2001-05-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.05" eventid="31" heat="2" lane="5">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="-1" lane="5" heat="2" heatid="20031" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Cape Verde" shortname="CPV" code="CPV" nation="CPV" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154801" lastname="PINA" firstname="Troy" gender="M" birthdate="1999-02-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.28" eventid="5" heat="3" lane="7">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="23" heat="1" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="59" lane="7" heat="3" heatid="30005" swimtime="00:00:26.90" reactiontime="+61" points="528">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:26.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="36" lane="3" heat="1" heatid="10023" swimtime="00:01:04.65" reactiontime="+62" points="442">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.50" />
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="75" swimtime="00:00:48.69" />
                    <SPLIT distance="100" swimtime="00:01:04.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154802" lastname="PINA" firstname="Jayla" gender="F" birthdate="2004-07-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.80" eventid="15" heat="2" lane="1">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="41" lane="1" heat="2" heatid="20015" swimtime="00:01:12.72" reactiontime="+67" points="630">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.37" />
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                    <SPLIT distance="75" swimtime="00:00:52.35" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="24" lane="1" heat="1" heatid="10022" swimtime="00:01:05.18" reactiontime="+70" points="651">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="75" swimtime="00:00:49.15" />
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Croatia" shortname="CRO" code="CRO" nation="CRO" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="125259" lastname="MILJENIC" firstname="Nikola" gender="M" birthdate="1998-05-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.23" eventid="39" heat="6" lane="7">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.37" eventid="14" heat="8" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.20" eventid="5" heat="6" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.14" eventid="31" heat="7" lane="8">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.54" eventid="23" heat="5" lane="8">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="20" lane="7" heat="6" heatid="60039" swimtime="00:00:51.16" reactiontime="+74" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.70" />
                    <SPLIT distance="50" swimtime="00:00:23.48" />
                    <SPLIT distance="75" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:00:51.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="30" lane="5" heat="8" heatid="80014" swimtime="00:00:47.51" reactiontime="+68" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.66" />
                    <SPLIT distance="50" swimtime="00:00:22.53" />
                    <SPLIT distance="75" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:00:47.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="26" lane="5" heat="6" heatid="60005" swimtime="00:00:22.90" reactiontime="+69" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.42" />
                    <SPLIT distance="50" swimtime="00:00:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="23" lane="8" heat="7" heatid="70031" swimtime="00:00:21.37" reactiontime="+71" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.32" />
                    <SPLIT distance="50" swimtime="00:00:21.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="20" lane="8" heat="5" heatid="50023" swimtime="00:00:52.85" reactiontime="+70" points="810">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.69" />
                    <SPLIT distance="50" swimtime="00:00:24.66" />
                    <SPLIT distance="75" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:00:52.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="115363" lastname="KAJTAZ" firstname="Amina" gender="F" birthdate="1996-12-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.98" eventid="38" heat="3" lane="1">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.63" eventid="20" heat="2" lane="2">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="18" lane="1" heat="3" heatid="30038" swimtime="00:00:57.88" reactiontime="+67" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="75" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:00:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="11" lane="2" heat="2" heatid="20020" swimtime="00:02:06.90" reactiontime="+54" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                    <SPLIT distance="75" swimtime="00:00:45.03" />
                    <SPLIT distance="100" swimtime="00:01:01.45" />
                    <SPLIT distance="125" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:01:33.57" />
                    <SPLIT distance="175" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:06.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182848" lastname="BOŠNJAK" firstname="Klara" gender="F" birthdate="2004-05-27">
              <ENTRIES>
                <ENTRY entrytime="00:08:47.11" eventid="12" heat="1" lane="3">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:16:51.57" eventid="33" heat="2" lane="1">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="17" lane="3" heat="1" heatid="10012" swimtime="00:08:49.67" reactiontime="+86" points="741">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="75" swimtime="00:00:46.73" />
                    <SPLIT distance="100" swimtime="00:01:03.12" />
                    <SPLIT distance="125" swimtime="00:01:19.60" />
                    <SPLIT distance="150" swimtime="00:01:36.01" />
                    <SPLIT distance="175" swimtime="00:01:52.62" />
                    <SPLIT distance="200" swimtime="00:02:09.18" />
                    <SPLIT distance="225" swimtime="00:02:25.78" />
                    <SPLIT distance="250" swimtime="00:02:42.26" />
                    <SPLIT distance="275" swimtime="00:02:58.89" />
                    <SPLIT distance="300" swimtime="00:03:15.56" />
                    <SPLIT distance="325" swimtime="00:03:32.25" />
                    <SPLIT distance="350" swimtime="00:03:48.98" />
                    <SPLIT distance="375" swimtime="00:04:05.75" />
                    <SPLIT distance="400" swimtime="00:04:22.59" />
                    <SPLIT distance="425" swimtime="00:04:39.35" />
                    <SPLIT distance="450" swimtime="00:04:56.14" />
                    <SPLIT distance="475" swimtime="00:05:13.03" />
                    <SPLIT distance="500" swimtime="00:05:29.88" />
                    <SPLIT distance="525" swimtime="00:05:46.50" />
                    <SPLIT distance="550" swimtime="00:06:03.34" />
                    <SPLIT distance="575" swimtime="00:06:20.08" />
                    <SPLIT distance="600" swimtime="00:06:36.87" />
                    <SPLIT distance="625" swimtime="00:06:53.43" />
                    <SPLIT distance="650" swimtime="00:07:10.15" />
                    <SPLIT distance="675" swimtime="00:07:26.86" />
                    <SPLIT distance="700" swimtime="00:07:43.71" />
                    <SPLIT distance="725" swimtime="00:08:00.38" />
                    <SPLIT distance="750" swimtime="00:08:16.88" />
                    <SPLIT distance="775" swimtime="00:08:33.67" />
                    <SPLIT distance="800" swimtime="00:08:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="14" lane="1" heat="2" heatid="20033" swimtime="00:16:51.02" reactiontime="+85" points="748">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.51" />
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="75" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:03.35" />
                    <SPLIT distance="125" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:01:36.56" />
                    <SPLIT distance="175" swimtime="00:01:53.35" />
                    <SPLIT distance="200" swimtime="00:02:10.19" />
                    <SPLIT distance="225" swimtime="00:02:27.04" />
                    <SPLIT distance="250" swimtime="00:02:43.80" />
                    <SPLIT distance="275" swimtime="00:03:00.53" />
                    <SPLIT distance="300" swimtime="00:03:17.45" />
                    <SPLIT distance="325" swimtime="00:03:34.31" />
                    <SPLIT distance="350" swimtime="00:03:51.19" />
                    <SPLIT distance="375" swimtime="00:04:08.01" />
                    <SPLIT distance="400" swimtime="00:04:25.05" />
                    <SPLIT distance="425" swimtime="00:04:41.97" />
                    <SPLIT distance="450" swimtime="00:04:59.01" />
                    <SPLIT distance="475" swimtime="00:05:15.98" />
                    <SPLIT distance="500" swimtime="00:05:33.10" />
                    <SPLIT distance="525" swimtime="00:05:50.14" />
                    <SPLIT distance="550" swimtime="00:06:07.11" />
                    <SPLIT distance="575" swimtime="00:06:24.24" />
                    <SPLIT distance="600" swimtime="00:06:41.19" />
                    <SPLIT distance="625" swimtime="00:06:58.15" />
                    <SPLIT distance="650" swimtime="00:07:15.18" />
                    <SPLIT distance="675" swimtime="00:07:32.21" />
                    <SPLIT distance="700" swimtime="00:07:49.27" />
                    <SPLIT distance="725" swimtime="00:08:06.19" />
                    <SPLIT distance="750" swimtime="00:08:23.26" />
                    <SPLIT distance="775" swimtime="00:08:40.27" />
                    <SPLIT distance="800" swimtime="00:08:57.20" />
                    <SPLIT distance="825" swimtime="00:09:14.19" />
                    <SPLIT distance="850" swimtime="00:09:31.16" />
                    <SPLIT distance="875" swimtime="00:09:48.09" />
                    <SPLIT distance="900" swimtime="00:10:05.13" />
                    <SPLIT distance="925" swimtime="00:10:22.31" />
                    <SPLIT distance="950" swimtime="00:10:39.41" />
                    <SPLIT distance="975" swimtime="00:10:56.49" />
                    <SPLIT distance="1000" swimtime="00:11:13.60" />
                    <SPLIT distance="1025" swimtime="00:11:30.71" />
                    <SPLIT distance="1050" swimtime="00:11:47.79" />
                    <SPLIT distance="1075" swimtime="00:12:04.70" />
                    <SPLIT distance="1100" swimtime="00:12:21.71" />
                    <SPLIT distance="1125" swimtime="00:12:38.39" />
                    <SPLIT distance="1150" swimtime="00:12:55.68" />
                    <SPLIT distance="1175" swimtime="00:13:12.67" />
                    <SPLIT distance="1200" swimtime="00:13:29.59" />
                    <SPLIT distance="1225" swimtime="00:13:46.41" />
                    <SPLIT distance="1250" swimtime="00:14:03.49" />
                    <SPLIT distance="1275" swimtime="00:14:20.27" />
                    <SPLIT distance="1300" swimtime="00:14:37.33" />
                    <SPLIT distance="1325" swimtime="00:14:54.27" />
                    <SPLIT distance="1350" swimtime="00:15:11.38" />
                    <SPLIT distance="1375" swimtime="00:15:28.14" />
                    <SPLIT distance="1400" swimtime="00:15:44.88" />
                    <SPLIT distance="1425" swimtime="00:16:01.50" />
                    <SPLIT distance="1450" swimtime="00:16:18.25" />
                    <SPLIT distance="1475" swimtime="00:16:34.90" />
                    <SPLIT distance="1500" swimtime="00:16:51.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Cuba" shortname="CUB" code="CUB" nation="CUB" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="101524" lastname="GAMEZ MATOS" firstname="Elisbet" gender="F" birthdate="1997-01-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.14" eventid="13" heat="6" lane="1">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.26" eventid="43" heat="4" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:04:09.08" eventid="1" heat="2" lane="2">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="34" lane="1" heat="6" heatid="60013" swimtime="00:00:54.87" reactiontime="+61" points="768">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:00:54.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="17" lane="7" heat="4" heatid="40043" swimtime="00:01:57.11" reactiontime="+62" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="75" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:00:57.73" />
                    <SPLIT distance="125" swimtime="00:01:12.61" />
                    <SPLIT distance="150" swimtime="00:01:27.58" />
                    <SPLIT distance="175" swimtime="00:01:42.70" />
                    <SPLIT distance="200" swimtime="00:01:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="18" lane="2" heat="2" heatid="20001" swimtime="00:04:11.66" reactiontime="+65" points="803">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="75" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:00:59.97" />
                    <SPLIT distance="125" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:31.32" />
                    <SPLIT distance="175" swimtime="00:01:47.19" />
                    <SPLIT distance="200" swimtime="00:02:03.27" />
                    <SPLIT distance="225" swimtime="00:02:19.28" />
                    <SPLIT distance="250" swimtime="00:02:35.42" />
                    <SPLIT distance="275" swimtime="00:02:51.55" />
                    <SPLIT distance="300" swimtime="00:03:07.64" />
                    <SPLIT distance="325" swimtime="00:03:23.62" />
                    <SPLIT distance="350" swimtime="00:03:39.94" />
                    <SPLIT distance="375" swimtime="00:03:56.02" />
                    <SPLIT distance="400" swimtime="00:04:11.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154025" lastname="FALCON JR." firstname="Rodolfo" gender="M" birthdate="2001-12-26">
              <ENTRIES>
                <ENTRY entrytime="00:08:24.45" eventid="42" heat="1" lane="1">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="142" place="20" lane="1" heat="1" heatid="10042" swimtime="00:08:11.47" reactiontime="+65" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="75" swimtime="00:00:42.78" />
                    <SPLIT distance="100" swimtime="00:00:57.94" />
                    <SPLIT distance="125" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:28.43" />
                    <SPLIT distance="175" swimtime="00:01:43.70" />
                    <SPLIT distance="200" swimtime="00:01:59.03" />
                    <SPLIT distance="225" swimtime="00:02:14.39" />
                    <SPLIT distance="250" swimtime="00:02:29.93" />
                    <SPLIT distance="275" swimtime="00:02:45.43" />
                    <SPLIT distance="300" swimtime="00:03:01.02" />
                    <SPLIT distance="325" swimtime="00:03:16.43" />
                    <SPLIT distance="350" swimtime="00:03:31.73" />
                    <SPLIT distance="375" swimtime="00:03:47.26" />
                    <SPLIT distance="400" swimtime="00:04:02.55" />
                    <SPLIT distance="425" swimtime="00:04:17.97" />
                    <SPLIT distance="450" swimtime="00:04:33.27" />
                    <SPLIT distance="475" swimtime="00:04:48.75" />
                    <SPLIT distance="500" swimtime="00:05:04.34" />
                    <SPLIT distance="525" swimtime="00:05:19.90" />
                    <SPLIT distance="550" swimtime="00:05:35.53" />
                    <SPLIT distance="575" swimtime="00:05:51.22" />
                    <SPLIT distance="600" swimtime="00:06:06.97" />
                    <SPLIT distance="625" swimtime="00:06:22.70" />
                    <SPLIT distance="650" swimtime="00:06:38.34" />
                    <SPLIT distance="675" swimtime="00:06:54.13" />
                    <SPLIT distance="700" swimtime="00:07:09.72" />
                    <SPLIT distance="725" swimtime="00:07:25.59" />
                    <SPLIT distance="750" swimtime="00:07:41.31" />
                    <SPLIT distance="775" swimtime="00:07:56.80" />
                    <SPLIT distance="800" swimtime="00:08:11.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Cyprus" shortname="CYP" code="CYP" nation="CYP" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="214214" lastname="HADJILOIZOU" firstname="Anna" gender="F" birthdate="2004-10-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.48" eventid="13" heat="5" lane="8">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.44" eventid="30" heat="5" lane="2">
                  <MEETINFO date="2022-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="29" lane="8" heat="5" heatid="50013" swimtime="00:00:54.52" reactiontime="+65" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                    <SPLIT distance="75" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:00:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="20" lane="2" heat="5" heatid="50030" swimtime="00:00:24.93" reactiontime="+63" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.16" />
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Czech Republic" shortname="CZE" code="CZE" nation="CZE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="110204" lastname="FRANTA" firstname="Tomas" gender="M" birthdate="1998-04-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.59" eventid="3" heat="5" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.36" eventid="19" heat="5" lane="2">
                  <MEETINFO date="2022-10-15" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="12" lane="6" heat="5" heatid="50003" swimtime="00:00:50.60" reactiontime="+61" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:24.53" />
                    <SPLIT distance="75" swimtime="00:00:37.49" />
                    <SPLIT distance="100" swimtime="00:00:50.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="11" lane="7" heat="1" heatid="10203" swimtime="00:00:50.39" reactiontime="+64" points="882">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:24.11" />
                    <SPLIT distance="75" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:00:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="13" lane="2" heat="5" heatid="50019" swimtime="00:00:23.26" reactiontime="+59" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.34" />
                    <SPLIT distance="50" swimtime="00:00:23.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="-1" lane="1" heat="2" heatid="20219" swimtime="00:00:23.05" status="DSQ" reactiontime="+58" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191812" lastname="ZABOJNIK" firstname="Matej" gender="M" birthdate="2000-08-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.59" eventid="16" heat="8" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.67" eventid="29" heat="4" lane="6">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:26.96" eventid="41" heat="6" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="16" lane="8" heat="8" heatid="80016" swimtime="00:00:57.87" reactiontime="+74" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="75" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:00:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="14" lane="8" heat="1" heatid="10216" swimtime="00:00:57.94" reactiontime="+75" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                    <SPLIT distance="75" swimtime="00:00:42.31" />
                    <SPLIT distance="100" swimtime="00:00:57.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="9" lane="6" heat="4" heatid="40029" swimtime="00:02:04.57" reactiontime="+72" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.45" />
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="75" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:00:59.07" />
                    <SPLIT distance="125" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:31.35" />
                    <SPLIT distance="175" swimtime="00:01:47.89" />
                    <SPLIT distance="200" swimtime="00:02:04.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="30" lane="6" heat="6" heatid="60041" swimtime="00:00:27.16" reactiontime="+70" points="775">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.25" />
                    <SPLIT distance="50" swimtime="00:00:27.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101618" lastname="SEFL" firstname="Jan" gender="M" birthdate="1990-05-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.46" eventid="39" heat="8" lane="8">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.53" eventid="5" heat="6" lane="8">
                  <MEETINFO date="2022-04-10" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.23" eventid="23" heat="4" lane="1">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="12" lane="8" heat="8" heatid="80039" swimtime="00:00:50.44" reactiontime="+69" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.66" />
                    <SPLIT distance="50" swimtime="00:00:23.50" />
                    <SPLIT distance="75" swimtime="00:00:36.61" />
                    <SPLIT distance="100" swimtime="00:00:50.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="16" lane="7" heat="1" heatid="10239" swimtime="00:00:51.03" reactiontime="+71" points="820">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.74" />
                    <SPLIT distance="50" swimtime="00:00:23.62" />
                    <SPLIT distance="75" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:00:51.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="24" lane="8" heat="6" heatid="60005" swimtime="00:00:22.84" reactiontime="+70" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.38" />
                    <SPLIT distance="50" swimtime="00:00:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="26" lane="1" heat="4" heatid="40023" swimtime="00:00:54.11" reactiontime="+67" points="755">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.60" />
                    <SPLIT distance="50" swimtime="00:00:24.28" />
                    <SPLIT distance="75" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:00:54.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210501" lastname="GRACIK" firstname="Daniel" gender="M" birthdate="2004-10-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.39" eventid="14" heat="7" lane="6">
                  <MEETINFO date="2022-10-14" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.46" eventid="5" heat="6" lane="6">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="41" lane="6" heat="7" heatid="70014" swimtime="00:00:48.14" reactiontime="+70" points="808">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.80" />
                    <SPLIT distance="50" swimtime="00:00:22.83" />
                    <SPLIT distance="75" swimtime="00:00:35.43" />
                    <SPLIT distance="100" swimtime="00:00:48.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="42" lane="6" heat="6" heatid="60005" swimtime="00:00:23.36" reactiontime="+72" points="807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.77" />
                    <SPLIT distance="50" swimtime="00:00:23.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149322" lastname="GEMOV" firstname="Ondřej" gender="M" birthdate="1999-06-12">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.69" eventid="21" heat="4" lane="7">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:07:50.16" eventid="42" heat="2" lane="1">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="21" place="15" lane="7" heat="4" heatid="40021" swimtime="00:01:52.92" reactiontime="+64" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:24.97" />
                    <SPLIT distance="75" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:00:53.33" />
                    <SPLIT distance="125" swimtime="00:01:07.88" />
                    <SPLIT distance="150" swimtime="00:01:22.71" />
                    <SPLIT distance="175" swimtime="00:01:37.75" />
                    <SPLIT distance="200" swimtime="00:01:52.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="10" lane="1" heat="2" heatid="20042" swimtime="00:07:42.70" reactiontime="+62" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:25.41" />
                    <SPLIT distance="75" swimtime="00:00:39.25" />
                    <SPLIT distance="100" swimtime="00:00:53.28" />
                    <SPLIT distance="125" swimtime="00:01:07.44" />
                    <SPLIT distance="150" swimtime="00:01:21.56" />
                    <SPLIT distance="175" swimtime="00:01:35.78" />
                    <SPLIT distance="200" swimtime="00:01:50.10" />
                    <SPLIT distance="225" swimtime="00:02:04.42" />
                    <SPLIT distance="250" swimtime="00:02:18.87" />
                    <SPLIT distance="275" swimtime="00:02:33.25" />
                    <SPLIT distance="300" swimtime="00:02:47.73" />
                    <SPLIT distance="325" swimtime="00:03:02.33" />
                    <SPLIT distance="350" swimtime="00:03:16.97" />
                    <SPLIT distance="375" swimtime="00:03:31.48" />
                    <SPLIT distance="400" swimtime="00:03:46.14" />
                    <SPLIT distance="425" swimtime="00:04:00.81" />
                    <SPLIT distance="450" swimtime="00:04:15.53" />
                    <SPLIT distance="475" swimtime="00:04:30.23" />
                    <SPLIT distance="500" swimtime="00:04:45.01" />
                    <SPLIT distance="525" swimtime="00:04:59.87" />
                    <SPLIT distance="550" swimtime="00:05:14.77" />
                    <SPLIT distance="575" swimtime="00:05:29.61" />
                    <SPLIT distance="600" swimtime="00:05:44.50" />
                    <SPLIT distance="625" swimtime="00:05:59.18" />
                    <SPLIT distance="650" swimtime="00:06:13.99" />
                    <SPLIT distance="675" swimtime="00:06:28.80" />
                    <SPLIT distance="700" swimtime="00:06:43.58" />
                    <SPLIT distance="725" swimtime="00:06:58.35" />
                    <SPLIT distance="750" swimtime="00:07:13.26" />
                    <SPLIT distance="775" swimtime="00:07:28.24" />
                    <SPLIT distance="800" swimtime="00:07:42.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214159" lastname="BURSA" firstname="Jakub" gender="M" birthdate="2003-01-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.72" eventid="7" heat="3" lane="8">
                  <MEETINFO date="2022-10-15" />
                </ENTRY>
                <ENTRY entrytime="00:04:09.06" eventid="37" heat="2" lane="1">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="25" lane="8" heat="3" heatid="30007" swimtime="00:01:58.01" reactiontime="+73" points="801">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:25.94" />
                    <SPLIT distance="75" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:00:55.87" />
                    <SPLIT distance="125" swimtime="00:01:12.39" />
                    <SPLIT distance="150" swimtime="00:01:29.58" />
                    <SPLIT distance="175" swimtime="00:01:44.55" />
                    <SPLIT distance="200" swimtime="00:01:58.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="14" lane="1" heat="2" heatid="20037" swimtime="00:04:10.28" reactiontime="+70" points="825">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.77" />
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                    <SPLIT distance="75" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:00:56.74" />
                    <SPLIT distance="125" swimtime="00:01:13.12" />
                    <SPLIT distance="150" swimtime="00:01:28.92" />
                    <SPLIT distance="175" swimtime="00:01:44.79" />
                    <SPLIT distance="200" swimtime="00:02:00.28" />
                    <SPLIT distance="225" swimtime="00:02:17.25" />
                    <SPLIT distance="250" swimtime="00:02:34.92" />
                    <SPLIT distance="275" swimtime="00:02:53.02" />
                    <SPLIT distance="300" swimtime="00:03:11.26" />
                    <SPLIT distance="325" swimtime="00:03:26.62" />
                    <SPLIT distance="350" swimtime="00:03:41.26" />
                    <SPLIT distance="375" swimtime="00:03:55.93" />
                    <SPLIT distance="400" swimtime="00:04:10.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101892" lastname="KUBOVA" firstname="Simona" gender="F" birthdate="1991-08-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.68" eventid="2" heat="4" lane="3">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.68" eventid="45" heat="5" lane="8">
                  <MEETINFO date="2021-09-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.38" eventid="18" heat="7" lane="2">
                  <MEETINFO date="2021-12-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="6" lane="3" heat="4" heatid="40002" swimtime="00:00:56.76" reactiontime="+57" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="75" swimtime="00:00:41.88" />
                    <SPLIT distance="100" swimtime="00:00:56.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="11" lane="3" heat="1" heatid="10202" swimtime="00:00:56.80" reactiontime="+60" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.36" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:41.95" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="19" lane="8" heat="5" heatid="50045" swimtime="00:02:06.19" reactiontime="+57" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="75" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:02.35" />
                    <SPLIT distance="125" swimtime="00:01:18.30" />
                    <SPLIT distance="150" swimtime="00:01:34.15" />
                    <SPLIT distance="175" swimtime="00:01:50.28" />
                    <SPLIT distance="200" swimtime="00:02:06.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="9" lane="2" heat="7" heatid="70018" swimtime="00:00:26.17" reactiontime="+56" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="12" lane="2" heat="2" heatid="20218" swimtime="00:00:26.32" reactiontime="+57" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121008" lastname="HORSKA" firstname="Kristyna" gender="F" birthdate="1997-09-30">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.60" eventid="15" heat="4" lane="2">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.89" eventid="28" heat="5" lane="3">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.85" eventid="6" heat="3" lane="2">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:01:00.31" eventid="22" heat="4" lane="2">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="29" lane="2" heat="4" heatid="40015" swimtime="00:01:06.57" reactiontime="+69" points="822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="75" swimtime="00:00:48.77" />
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="13" lane="3" heat="5" heatid="50028" swimtime="00:02:21.22" reactiontime="+71" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="75" swimtime="00:00:49.72" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="125" swimtime="00:01:25.74" />
                    <SPLIT distance="150" swimtime="00:01:43.96" />
                    <SPLIT distance="175" swimtime="00:02:02.31" />
                    <SPLIT distance="200" swimtime="00:02:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="20" lane="2" heat="3" heatid="30006" swimtime="00:02:10.46" reactiontime="+72" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.61" />
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                    <SPLIT distance="75" swimtime="00:00:45.75" />
                    <SPLIT distance="100" swimtime="00:01:02.22" />
                    <SPLIT distance="125" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:01:38.91" />
                    <SPLIT distance="175" swimtime="00:01:55.45" />
                    <SPLIT distance="200" swimtime="00:02:10.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="-1" lane="2" heat="4" heatid="40022" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120699" lastname="JANICKOVA" firstname="Barbora" gender="F" birthdate="2000-05-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.33" eventid="38" heat="2" lane="8">
                  <MEETINFO date="2021-10-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.75" eventid="13" heat="9" lane="8">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="21" lane="8" heat="2" heatid="20038" swimtime="00:00:58.65" reactiontime="+69" points="806">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                    <SPLIT distance="75" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:00:58.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="18" lane="8" heat="9" heatid="90013" swimtime="00:00:53.45" reactiontime="+68" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:25.62" />
                    <SPLIT distance="75" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:00:53.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="120507" lastname="SEEMANOVA" firstname="Barbora" gender="F" birthdate="2000-04-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.71" eventid="13" heat="7" lane="5">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.23" eventid="43" heat="5" lane="3">
                  <MEETINFO date="2021-11-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.23" eventid="4" heat="5" lane="1">
                  <MEETINFO date="2022-10-15" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.26" eventid="30" heat="8" lane="7">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="7" lane="5" heat="7" heatid="70013" swimtime="00:00:52.54" reactiontime="+61" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:25.22" />
                    <SPLIT distance="75" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="12" lane="6" heat="2" heatid="20213" swimtime="00:00:52.59" reactiontime="+62" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:25.10" />
                    <SPLIT distance="75" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:00:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="143" place="5" lane="6" heat="1" heatid="10143" swimtime="00:01:52.66" reactiontime="+61" points="938">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="75" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:00:54.49" />
                    <SPLIT distance="125" swimtime="00:01:08.97" />
                    <SPLIT distance="150" swimtime="00:01:23.57" />
                    <SPLIT distance="175" swimtime="00:01:38.29" />
                    <SPLIT distance="200" swimtime="00:01:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="4" lane="3" heat="5" heatid="50043" swimtime="00:01:53.67" reactiontime="+61" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.45" />
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                    <SPLIT distance="75" swimtime="00:00:41.04" />
                    <SPLIT distance="100" swimtime="00:00:55.74" />
                    <SPLIT distance="125" swimtime="00:01:10.35" />
                    <SPLIT distance="150" swimtime="00:01:24.93" />
                    <SPLIT distance="175" swimtime="00:01:39.54" />
                    <SPLIT distance="200" swimtime="00:01:53.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="21" lane="1" heat="5" heatid="50004" swimtime="00:00:26.09" reactiontime="+64" points="815">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="11" lane="7" heat="8" heatid="80030" swimtime="00:00:24.24" reactiontime="+63" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:24.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="13" lane="7" heat="2" heatid="20230" swimtime="00:00:24.25" reactiontime="+60" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:24.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Czech Republic">
              <RESULTS>
                <RESULT eventid="148" place="8" lane="8" heat="1" swimtime="00:03:26.37" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.54" />
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="75" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:00:50.48" />
                    <SPLIT distance="125" swimtime="00:01:02.25" />
                    <SPLIT distance="150" swimtime="00:01:17.08" />
                    <SPLIT distance="175" swimtime="00:01:32.13" />
                    <SPLIT distance="200" swimtime="00:01:47.97" />
                    <SPLIT distance="225" swimtime="00:01:58.30" />
                    <SPLIT distance="250" swimtime="00:02:11.18" />
                    <SPLIT distance="275" swimtime="00:02:24.63" />
                    <SPLIT distance="300" swimtime="00:02:38.75" />
                    <SPLIT distance="325" swimtime="00:02:48.94" />
                    <SPLIT distance="350" swimtime="00:03:01.27" />
                    <SPLIT distance="375" swimtime="00:03:13.74" />
                    <SPLIT distance="400" swimtime="00:03:26.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="110204" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="191812" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="101618" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="210501" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="8" lane="5" heat="1" swimtime="00:03:26.18" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                    <SPLIT distance="75" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:00:50.42" />
                    <SPLIT distance="125" swimtime="00:01:02.36" />
                    <SPLIT distance="150" swimtime="00:01:17.04" />
                    <SPLIT distance="175" swimtime="00:01:32.18" />
                    <SPLIT distance="200" swimtime="00:01:47.84" />
                    <SPLIT distance="225" swimtime="00:01:58.07" />
                    <SPLIT distance="250" swimtime="00:02:10.90" />
                    <SPLIT distance="275" swimtime="00:02:24.26" />
                    <SPLIT distance="300" swimtime="00:02:38.32" />
                    <SPLIT distance="325" swimtime="00:02:48.74" />
                    <SPLIT distance="350" swimtime="00:03:00.71" />
                    <SPLIT distance="375" swimtime="00:03:13.51" />
                    <SPLIT distance="400" swimtime="00:03:26.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="110204" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="191812" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="101618" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="210501" reactiontime="+45" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Czech Republic">
              <RESULTS>
                <RESULT eventid="134" place="8" lane="8" heat="1" swimtime="00:01:46.40" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="75" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:00:56.90" />
                    <SPLIT distance="125" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:22.33" />
                    <SPLIT distance="175" swimtime="00:01:33.83" />
                    <SPLIT distance="200" swimtime="00:01:46.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101892" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="121008" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="120507" reactiontime="+33" />
                    <RELAYPOSITION number="4" athleteid="120699" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="8" lane="7" heat="1" swimtime="00:01:46.73" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                    <SPLIT distance="75" swimtime="00:00:40.17" />
                    <SPLIT distance="100" swimtime="00:00:57.13" />
                    <SPLIT distance="125" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:22.65" />
                    <SPLIT distance="175" swimtime="00:01:34.16" />
                    <SPLIT distance="200" swimtime="00:01:46.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101892" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="121008" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="120507" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="120699" reactiontime="+12" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Denmark" shortname="DEN" code="DEN" nation="DEN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="181160" lastname="BLOMSTERBERG" firstname="Thea" gender="F" birthdate="2002-01-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.54" eventid="15" heat="6" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.96" eventid="28" heat="3" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="11" lane="8" heat="6" heatid="60015" swimtime="00:01:04.74" reactiontime="+67" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="75" swimtime="00:00:47.74" />
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="13" lane="7" heat="2" heatid="20215" swimtime="00:01:05.22" reactiontime="+72" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="75" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="128" place="7" lane="1" heat="1" heatid="10128" swimtime="00:02:20.14" reactiontime="+73" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="75" swimtime="00:00:49.04" />
                    <SPLIT distance="100" swimtime="00:01:06.79" />
                    <SPLIT distance="125" swimtime="00:01:24.73" />
                    <SPLIT distance="150" swimtime="00:01:42.94" />
                    <SPLIT distance="175" swimtime="00:02:01.18" />
                    <SPLIT distance="200" swimtime="00:02:20.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="7" lane="3" heat="3" heatid="30028" swimtime="00:02:19.88" reactiontime="+69" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.94" />
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="75" swimtime="00:00:49.46" />
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="125" swimtime="00:01:25.25" />
                    <SPLIT distance="150" swimtime="00:01:43.47" />
                    <SPLIT distance="175" swimtime="00:02:01.57" />
                    <SPLIT distance="200" swimtime="00:02:19.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191642" lastname="BACH" firstname="Helena" gender="F" birthdate="2000-06-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.73" eventid="38" heat="3" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.02" eventid="20" heat="2" lane="5">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.66" eventid="43" heat="5" lane="1">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="00:04:04.11" eventid="1" heat="3" lane="1">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="11" lane="7" heat="3" heatid="30038" swimtime="00:00:57.15" reactiontime="+78" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:00:57.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="13" lane="7" heat="2" heatid="20238" swimtime="00:00:57.21" reactiontime="+78" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:00:57.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="120" place="4" lane="3" heat="1" heatid="10120" swimtime="00:02:04.41" reactiontime="+76" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="75" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:00.14" />
                    <SPLIT distance="125" swimtime="00:01:15.93" />
                    <SPLIT distance="150" swimtime="00:01:32.13" />
                    <SPLIT distance="175" swimtime="00:01:48.16" />
                    <SPLIT distance="200" swimtime="00:02:04.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="3" lane="5" heat="2" heatid="20020" swimtime="00:02:05.09" reactiontime="+78" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.32" />
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="75" swimtime="00:00:44.73" />
                    <SPLIT distance="100" swimtime="00:01:00.62" />
                    <SPLIT distance="125" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:32.64" />
                    <SPLIT distance="175" swimtime="00:01:48.82" />
                    <SPLIT distance="200" swimtime="00:02:05.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="12" lane="1" heat="5" heatid="50043" swimtime="00:01:55.79" reactiontime="+78" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                    <SPLIT distance="75" swimtime="00:00:41.89" />
                    <SPLIT distance="100" swimtime="00:00:56.50" />
                    <SPLIT distance="125" swimtime="00:01:11.14" />
                    <SPLIT distance="150" swimtime="00:01:26.06" />
                    <SPLIT distance="175" swimtime="00:01:41.20" />
                    <SPLIT distance="200" swimtime="00:01:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="10" lane="1" heat="3" heatid="30001" swimtime="00:04:03.59" reactiontime="+76" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.64" />
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="75" swimtime="00:00:43.81" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="125" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:01:29.52" />
                    <SPLIT distance="175" swimtime="00:01:44.79" />
                    <SPLIT distance="200" swimtime="00:02:00.18" />
                    <SPLIT distance="225" swimtime="00:02:15.41" />
                    <SPLIT distance="250" swimtime="00:02:30.82" />
                    <SPLIT distance="275" swimtime="00:02:46.16" />
                    <SPLIT distance="300" swimtime="00:03:01.75" />
                    <SPLIT distance="325" swimtime="00:03:17.24" />
                    <SPLIT distance="350" swimtime="00:03:32.74" />
                    <SPLIT distance="375" swimtime="00:03:48.49" />
                    <SPLIT distance="400" swimtime="00:04:03.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106983" lastname="JENSEN" firstname="Julie Kepp" gender="F" birthdate="2000-01-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.25" eventid="18" heat="7" lane="6">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.31" eventid="4" heat="5" lane="6">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.03" eventid="30" heat="8" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="118" place="7" lane="1" heat="1" heatid="10118" swimtime="00:00:26.14" reactiontime="+59" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="1" lane="6" heat="7" heatid="70018" swimtime="00:00:25.85" reactiontime="+55" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="7" lane="4" heat="2" heatid="20218" swimtime="00:00:26.02" reactiontime="+57" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.69" />
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="14" lane="6" heat="5" heatid="50004" swimtime="00:00:25.51" reactiontime="+64" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="14" lane="1" heat="1" heatid="10204" swimtime="00:00:25.56" reactiontime="+64" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="4" lane="2" heat="1" heatid="10130" swimtime="00:00:23.71" reactiontime="+63" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="3" lane="2" heat="8" heatid="80030" swimtime="00:00:23.79" reactiontime="+60" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="5" lane="5" heat="2" heatid="20230" swimtime="00:00:23.93" reactiontime="+63" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:23.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Dominican Rep." shortname="DOM" code="DOM" nation="DOM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="108183" lastname="DOMINGUEZ RAMOS" firstname="Josue" gender="M" birthdate="1996-11-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.44" eventid="16" heat="5" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.91" eventid="41" heat="6" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="38" lane="6" heat="5" heatid="50016" swimtime="00:00:59.73" reactiontime="+62" points="792">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                    <SPLIT distance="75" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:00:59.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="32" lane="5" heat="6" heatid="60041" swimtime="00:00:27.18" reactiontime="+60" points="773">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149544" lastname="GONZALEZ RAMIREZ" firstname="Denzel" gender="M" birthdate="2000-02-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.43" eventid="39" heat="3" lane="6">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:50.13" eventid="14" heat="6" lane="8">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="42" lane="6" heat="3" heatid="30039" swimtime="00:00:54.90" reactiontime="+59" points="659">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.19" />
                    <SPLIT distance="50" swimtime="00:00:24.96" />
                    <SPLIT distance="75" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:00:54.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="47" lane="8" heat="6" heatid="60014" swimtime="00:00:49.59" reactiontime="+61" points="739">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.04" />
                    <SPLIT distance="50" swimtime="00:00:23.27" />
                    <SPLIT distance="75" swimtime="00:00:36.31" />
                    <SPLIT distance="100" swimtime="00:00:49.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197991" lastname="JIMENEZ" firstname="Elizabeth" gender="F" birthdate="2006-02-06">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:03.29" eventid="2" heat="2" lane="3">
                  <MEETINFO date="2022-04-02" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.23" eventid="45" heat="2" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="35" lane="3" heat="2" heatid="20002" swimtime="00:01:01.44" reactiontime="+61" points="713">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.35" />
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="75" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="31" lane="1" heat="2" heatid="20045" swimtime="00:02:12.63" reactiontime="+62" points="721">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.50" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:46.51" />
                    <SPLIT distance="100" swimtime="00:01:03.56" />
                    <SPLIT distance="125" swimtime="00:01:20.51" />
                    <SPLIT distance="150" swimtime="00:01:37.85" />
                    <SPLIT distance="175" swimtime="00:01:55.46" />
                    <SPLIT distance="200" swimtime="00:02:12.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="152506" lastname="LARA" firstname="Krystal" gender="F" birthdate="1998-03-18">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:00.66" eventid="38" heat="1" lane="4">
                  <MEETINFO date="2022-07-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.65" eventid="20" heat="1" lane="5">
                  <MEETINFO date="2022-07-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="24" lane="4" heat="1" heatid="10038" swimtime="00:00:59.78" reactiontime="+51" points="761">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="75" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:00:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="18" lane="5" heat="1" heatid="10020" swimtime="00:02:11.43" reactiontime="+67" points="753">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.49" />
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="75" swimtime="00:00:45.75" />
                    <SPLIT distance="100" swimtime="00:01:02.52" />
                    <SPLIT distance="125" swimtime="00:01:19.55" />
                    <SPLIT distance="150" swimtime="00:01:36.57" />
                    <SPLIT distance="175" swimtime="00:01:54.14" />
                    <SPLIT distance="200" swimtime="00:02:11.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Dominican Republic">
              <RESULTS>
                <RESULT eventid="27" place="17" lane="6" heat="3" swimtime="00:01:37.25" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.90" />
                    <SPLIT distance="50" swimtime="00:00:22.95" />
                    <SPLIT distance="75" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:00:49.42" />
                    <SPLIT distance="125" swimtime="00:01:01.28" />
                    <SPLIT distance="150" swimtime="00:01:14.77" />
                    <SPLIT distance="175" swimtime="00:01:25.33" />
                    <SPLIT distance="200" swimtime="00:01:37.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="108183" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="197991" reactiontime="+37" />
                    <RELAYPOSITION number="3" athleteid="152506" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="149544" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Dominican Republic">
              <RESULTS>
                <RESULT eventid="11" place="20" lane="6" heat="3" swimtime="00:01:44.73" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.30" />
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                    <SPLIT distance="75" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:00:55.17" />
                    <SPLIT distance="125" swimtime="00:01:07.53" />
                    <SPLIT distance="150" swimtime="00:01:22.48" />
                    <SPLIT distance="175" swimtime="00:01:32.93" />
                    <SPLIT distance="200" swimtime="00:01:44.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197991" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="108183" reactiontime="+11" />
                    <RELAYPOSITION number="3" athleteid="152506" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="149544" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Ecuador" shortname="ECU" code="ECU" nation="ECU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="120206" lastname="PERIBONIO AVILA" firstname="Tomas" gender="M" birthdate="1996-01-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.39" eventid="7" heat="5" lane="8">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="22" lane="8" heat="5" heatid="50007" swimtime="00:01:57.32" reactiontime="+63" points="815">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:25.10" />
                    <SPLIT distance="75" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:00:54.79" />
                    <SPLIT distance="125" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:28.21" />
                    <SPLIT distance="175" swimtime="00:01:43.21" />
                    <SPLIT distance="200" swimtime="00:01:57.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149867" lastname="DELGADO" firstname="Anicka" gender="F" birthdate="2002-06-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.56" eventid="13" heat="5" lane="2">
                  <MEETINFO date="2021-07-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.12" eventid="4" heat="3" lane="4">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="25" lane="2" heat="5" heatid="50013" swimtime="00:00:54.19" reactiontime="+67" points="797">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.25" />
                    <SPLIT distance="50" swimtime="00:00:26.03" />
                    <SPLIT distance="75" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:00:54.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="20" lane="4" heat="3" heatid="30004" swimtime="00:00:26.04" reactiontime="+66" points="820">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.00" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Egypt" shortname="EGY" code="EGY" nation="EGY" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="121963" lastname="ELKAMASH" firstname="Youssef" gender="M" birthdate="1995-07-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.18" eventid="16" heat="4" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.90" eventid="41" heat="6" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="36" lane="6" heat="4" heatid="40016" swimtime="00:00:59.61" reactiontime="+68" points="797">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="75" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:00:59.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="34" lane="4" heat="6" heatid="60041" swimtime="00:00:27.28" reactiontime="+66" points="765">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.51" />
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183396" lastname="RAMADAN" firstname="Youssef" gender="M" birthdate="2002-07-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.50" eventid="39" heat="6" lane="5">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:46.98" eventid="14" heat="11" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.63" eventid="5" heat="9" lane="7">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="8" lane="8" heat="1" heatid="10139" swimtime="00:00:49.84" reactiontime="+60" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.62" />
                    <SPLIT distance="50" swimtime="00:00:22.98" />
                    <SPLIT distance="75" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:00:49.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="3" lane="5" heat="6" heatid="60039" swimtime="00:00:49.64" reactiontime="+60" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.86" />
                    <SPLIT distance="50" swimtime="00:00:23.42" />
                    <SPLIT distance="75" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:00:49.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="8" lane="5" heat="2" heatid="20239" swimtime="00:00:49.79" reactiontime="+58" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.73" />
                    <SPLIT distance="50" swimtime="00:00:23.41" />
                    <SPLIT distance="75" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:00:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="8" lane="1" heat="11" heatid="110014" swimtime="00:00:46.51" reactiontime="+60" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.30" />
                    <SPLIT distance="50" swimtime="00:00:21.96" />
                    <SPLIT distance="75" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:00:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="10" lane="6" heat="1" heatid="10214" swimtime="00:00:46.57" reactiontime="+60" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.65" />
                    <SPLIT distance="50" swimtime="00:00:22.28" />
                    <SPLIT distance="75" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="15" lane="7" heat="9" heatid="90005" swimtime="00:00:22.50" reactiontime="+60" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.45" />
                    <SPLIT distance="50" swimtime="00:00:22.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="10" lane="8" heat="2" heatid="20205" swimtime="00:00:22.32" reactiontime="+60" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:22.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110774" lastname="ELKAMASH" firstname="Marwan" gender="M" birthdate="1993-11-14">
              <ENTRIES>
                <ENTRY entrytime="00:14:35.93" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.94" eventid="24" heat="5" lane="8">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:07:45.09" eventid="42" heat="2" lane="5">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="11" lane="1" heat="5" heatid="30110" swimtime="00:14:53.57" reactiontime="+71" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                    <SPLIT distance="75" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:00:55.29" />
                    <SPLIT distance="125" swimtime="00:01:09.91" />
                    <SPLIT distance="150" swimtime="00:01:24.41" />
                    <SPLIT distance="175" swimtime="00:01:39.04" />
                    <SPLIT distance="200" swimtime="00:01:53.47" />
                    <SPLIT distance="225" swimtime="00:02:08.24" />
                    <SPLIT distance="250" swimtime="00:02:22.69" />
                    <SPLIT distance="275" swimtime="00:02:37.13" />
                    <SPLIT distance="300" swimtime="00:02:51.53" />
                    <SPLIT distance="325" swimtime="00:03:06.22" />
                    <SPLIT distance="350" swimtime="00:03:20.64" />
                    <SPLIT distance="375" swimtime="00:03:35.07" />
                    <SPLIT distance="400" swimtime="00:03:49.56" />
                    <SPLIT distance="425" swimtime="00:04:04.05" />
                    <SPLIT distance="450" swimtime="00:04:18.64" />
                    <SPLIT distance="475" swimtime="00:04:33.36" />
                    <SPLIT distance="500" swimtime="00:04:48.14" />
                    <SPLIT distance="525" swimtime="00:05:03.03" />
                    <SPLIT distance="550" swimtime="00:05:18.11" />
                    <SPLIT distance="575" swimtime="00:05:33.25" />
                    <SPLIT distance="600" swimtime="00:05:48.34" />
                    <SPLIT distance="625" swimtime="00:06:03.39" />
                    <SPLIT distance="650" swimtime="00:06:18.41" />
                    <SPLIT distance="675" swimtime="00:06:33.53" />
                    <SPLIT distance="700" swimtime="00:06:48.97" />
                    <SPLIT distance="725" swimtime="00:07:04.39" />
                    <SPLIT distance="750" swimtime="00:07:19.75" />
                    <SPLIT distance="775" swimtime="00:07:34.96" />
                    <SPLIT distance="800" swimtime="00:07:50.41" />
                    <SPLIT distance="825" swimtime="00:08:05.63" />
                    <SPLIT distance="850" swimtime="00:08:21.13" />
                    <SPLIT distance="875" swimtime="00:08:36.22" />
                    <SPLIT distance="900" swimtime="00:08:51.37" />
                    <SPLIT distance="925" swimtime="00:09:06.71" />
                    <SPLIT distance="950" swimtime="00:09:21.95" />
                    <SPLIT distance="975" swimtime="00:09:37.30" />
                    <SPLIT distance="1000" swimtime="00:09:52.42" />
                    <SPLIT distance="1025" swimtime="00:10:07.59" />
                    <SPLIT distance="1050" swimtime="00:10:22.81" />
                    <SPLIT distance="1075" swimtime="00:10:37.83" />
                    <SPLIT distance="1100" swimtime="00:10:53.20" />
                    <SPLIT distance="1125" swimtime="00:11:08.06" />
                    <SPLIT distance="1150" swimtime="00:11:23.41" />
                    <SPLIT distance="1175" swimtime="00:11:38.55" />
                    <SPLIT distance="1200" swimtime="00:11:53.54" />
                    <SPLIT distance="1225" swimtime="00:12:08.45" />
                    <SPLIT distance="1250" swimtime="00:12:23.61" />
                    <SPLIT distance="1275" swimtime="00:12:38.60" />
                    <SPLIT distance="1300" swimtime="00:12:53.93" />
                    <SPLIT distance="1325" swimtime="00:13:08.95" />
                    <SPLIT distance="1350" swimtime="00:13:24.24" />
                    <SPLIT distance="1375" swimtime="00:13:39.57" />
                    <SPLIT distance="1400" swimtime="00:13:54.84" />
                    <SPLIT distance="1425" swimtime="00:14:09.48" />
                    <SPLIT distance="1450" swimtime="00:14:24.55" />
                    <SPLIT distance="1475" swimtime="00:14:39.24" />
                    <SPLIT distance="1500" swimtime="00:14:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="-1" lane="8" heat="5" heatid="50024" swimtime="NT" status="DNS" />
                <RESULT eventid="142" place="7" lane="5" heat="2" heatid="20042" swimtime="00:07:36.01" reactiontime="+71" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                    <SPLIT distance="75" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:00:55.35" />
                    <SPLIT distance="125" swimtime="00:01:09.87" />
                    <SPLIT distance="150" swimtime="00:01:24.40" />
                    <SPLIT distance="175" swimtime="00:01:38.83" />
                    <SPLIT distance="200" swimtime="00:01:53.28" />
                    <SPLIT distance="225" swimtime="00:02:07.89" />
                    <SPLIT distance="250" swimtime="00:02:22.29" />
                    <SPLIT distance="275" swimtime="00:02:36.73" />
                    <SPLIT distance="300" swimtime="00:02:51.11" />
                    <SPLIT distance="325" swimtime="00:03:05.55" />
                    <SPLIT distance="350" swimtime="00:03:19.98" />
                    <SPLIT distance="375" swimtime="00:03:34.38" />
                    <SPLIT distance="400" swimtime="00:03:48.74" />
                    <SPLIT distance="425" swimtime="00:04:03.15" />
                    <SPLIT distance="450" swimtime="00:04:17.52" />
                    <SPLIT distance="475" swimtime="00:04:32.00" />
                    <SPLIT distance="500" swimtime="00:04:46.32" />
                    <SPLIT distance="525" swimtime="00:05:00.78" />
                    <SPLIT distance="550" swimtime="00:05:15.10" />
                    <SPLIT distance="575" swimtime="00:05:29.43" />
                    <SPLIT distance="600" swimtime="00:05:43.61" />
                    <SPLIT distance="625" swimtime="00:05:57.85" />
                    <SPLIT distance="650" swimtime="00:06:11.98" />
                    <SPLIT distance="675" swimtime="00:06:26.19" />
                    <SPLIT distance="700" swimtime="00:06:40.33" />
                    <SPLIT distance="725" swimtime="00:06:54.48" />
                    <SPLIT distance="750" swimtime="00:07:08.61" />
                    <SPLIT distance="775" swimtime="00:07:22.57" />
                    <SPLIT distance="800" swimtime="00:07:36.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150480" lastname="SAMEH" firstname="Abdelrahman" gender="M" birthdate="2000-03-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:22.76" eventid="5" heat="8" lane="8">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="33" lane="8" heat="8" heatid="80005" swimtime="00:00:23.11" reactiontime="+63" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.46" />
                    <SPLIT distance="50" swimtime="00:00:23.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121964" lastname="KHALAFALLA" firstname="Ali" gender="M" birthdate="1996-05-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:21.37" eventid="31" heat="11" lane="8">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="22" lane="8" heat="11" heatid="110031" swimtime="00:00:21.36" reactiontime="+61" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.22" />
                    <SPLIT distance="50" swimtime="00:00:21.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="El Salvador" shortname="ESA" code="ESA" nation="ESA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="210623" lastname="VENTURA" firstname="Xavier" gender="M" birthdate="2007-03-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.66" eventid="39" heat="3" lane="1">
                  <MEETINFO date="2022-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.67" eventid="21" heat="2" lane="8">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="47" lane="1" heat="3" heatid="30039" swimtime="00:00:56.38" reactiontime="+69" points="608">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                    <SPLIT distance="75" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:00:56.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="23" lane="8" heat="2" heatid="20021" swimtime="00:02:02.63" reactiontime="+71" points="687">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                    <SPLIT distance="75" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:00:58.73" />
                    <SPLIT distance="125" swimtime="00:01:14.60" />
                    <SPLIT distance="150" swimtime="00:01:30.68" />
                    <SPLIT distance="175" swimtime="00:01:46.48" />
                    <SPLIT distance="200" swimtime="00:02:02.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108069" lastname="MARQUEZ" firstname="Celina" gender="F" birthdate="1999-07-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.82" eventid="2" heat="3" lane="1">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.23" eventid="45" heat="2" lane="6">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="33" lane="1" heat="3" heatid="30002" swimtime="00:01:01.08" reactiontime="+55" points="725">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="75" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:01:01.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="32" lane="6" heat="2" heatid="20045" swimtime="00:02:13.61" reactiontime="+55" points="705">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.99" />
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="75" swimtime="00:00:48.09" />
                    <SPLIT distance="100" swimtime="00:01:05.02" />
                    <SPLIT distance="125" swimtime="00:01:22.05" />
                    <SPLIT distance="150" swimtime="00:01:39.15" />
                    <SPLIT distance="175" swimtime="00:01:56.76" />
                    <SPLIT distance="200" swimtime="00:02:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Spain" shortname="ESP" code="ESP" nation="ESP" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154214" lastname="COLL MARTI" firstname="Carles" gender="M" birthdate="2001-10-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.56" eventid="16" heat="5" lane="7">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.17" eventid="29" heat="4" lane="7">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.31" eventid="7" heat="3" lane="2">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:52.36" eventid="23" heat="4" lane="2">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="-1" lane="7" heat="5" heatid="50016" swimtime="NT" status="DNS" />
                <RESULT eventid="29" place="-1" lane="7" heat="4" heatid="40029" swimtime="NT" status="DNS" />
                <RESULT eventid="7" place="13" lane="2" heat="3" heatid="30007" swimtime="00:01:54.03" reactiontime="+63" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.30" />
                    <SPLIT distance="50" swimtime="00:00:25.15" />
                    <SPLIT distance="75" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:00:53.36" />
                    <SPLIT distance="125" swimtime="00:01:09.17" />
                    <SPLIT distance="150" swimtime="00:01:25.67" />
                    <SPLIT distance="175" swimtime="00:01:40.38" />
                    <SPLIT distance="200" swimtime="00:01:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="8" lane="8" heat="1" heatid="10123" swimtime="00:00:52.36" reactiontime="+61" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.67" />
                    <SPLIT distance="50" swimtime="00:00:23.75" />
                    <SPLIT distance="75" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="9" lane="2" heat="4" heatid="40023" swimtime="00:00:52.32" reactiontime="+62" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.87" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                    <SPLIT distance="75" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="8" lane="2" heat="2" heatid="20223" swimtime="00:00:51.97" reactiontime="+60" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.59" />
                    <SPLIT distance="50" swimtime="00:00:23.53" />
                    <SPLIT distance="75" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:00:51.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182683" lastname="MOLLA YANES" firstname="Mario" gender="M" birthdate="2002-04-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.42" eventid="39" heat="5" lane="2">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.54" eventid="5" heat="5" lane="4">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="17" lane="2" heat="5" heatid="50039" swimtime="00:00:50.67" reactiontime="+64" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.42" />
                    <SPLIT distance="75" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:00:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="23" lane="4" heat="5" heatid="50005" swimtime="00:00:22.83" reactiontime="+63" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.43" />
                    <SPLIT distance="50" swimtime="00:00:22.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154217" lastname="DE CELIS MONTALBAN" firstname="Sergio" gender="M" birthdate="2000-01-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.41" eventid="14" heat="7" lane="1">
                  <MEETINFO date="2022-08-14" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.97" eventid="31" heat="7" lane="2">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="12" lane="1" heat="7" heatid="70014" swimtime="00:00:46.80" reactiontime="+65" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.52" />
                    <SPLIT distance="75" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:00:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="11" lane="7" heat="1" heatid="10214" swimtime="00:00:46.60" reactiontime="+67" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.74" />
                    <SPLIT distance="50" swimtime="00:00:22.63" />
                    <SPLIT distance="75" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:00:46.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="-1" lane="2" heat="7" heatid="70031" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201563" lastname="GARACH BENITO" firstname="Carlos" gender="M" birthdate="2004-07-25">
              <ENTRIES>
                <ENTRY entrytime="00:14:45.16" eventid="10" heat="2" lane="3">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="00:07:52.73" eventid="42" heat="1" lane="5">
                  <MEETINFO date="2022-09-01" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="14" lane="3" heat="2" heatid="20010" swimtime="00:14:59.37" reactiontime="+68" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                    <SPLIT distance="75" swimtime="00:00:40.26" />
                    <SPLIT distance="100" swimtime="00:00:54.53" />
                    <SPLIT distance="125" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:23.58" />
                    <SPLIT distance="175" swimtime="00:01:38.09" />
                    <SPLIT distance="200" swimtime="00:01:52.70" />
                    <SPLIT distance="225" swimtime="00:02:07.18" />
                    <SPLIT distance="250" swimtime="00:02:21.80" />
                    <SPLIT distance="275" swimtime="00:02:36.33" />
                    <SPLIT distance="300" swimtime="00:02:51.08" />
                    <SPLIT distance="325" swimtime="00:03:05.80" />
                    <SPLIT distance="350" swimtime="00:03:20.71" />
                    <SPLIT distance="375" swimtime="00:03:35.64" />
                    <SPLIT distance="400" swimtime="00:03:50.72" />
                    <SPLIT distance="425" swimtime="00:04:05.66" />
                    <SPLIT distance="450" swimtime="00:04:20.65" />
                    <SPLIT distance="475" swimtime="00:04:35.59" />
                    <SPLIT distance="500" swimtime="00:04:50.66" />
                    <SPLIT distance="525" swimtime="00:05:05.66" />
                    <SPLIT distance="550" swimtime="00:05:20.83" />
                    <SPLIT distance="575" swimtime="00:05:35.93" />
                    <SPLIT distance="600" swimtime="00:05:51.13" />
                    <SPLIT distance="625" swimtime="00:06:06.21" />
                    <SPLIT distance="650" swimtime="00:06:21.56" />
                    <SPLIT distance="675" swimtime="00:06:36.79" />
                    <SPLIT distance="700" swimtime="00:06:52.09" />
                    <SPLIT distance="725" swimtime="00:07:07.29" />
                    <SPLIT distance="750" swimtime="00:07:22.52" />
                    <SPLIT distance="775" swimtime="00:07:37.79" />
                    <SPLIT distance="800" swimtime="00:07:53.07" />
                    <SPLIT distance="825" swimtime="00:08:08.38" />
                    <SPLIT distance="850" swimtime="00:08:23.73" />
                    <SPLIT distance="875" swimtime="00:08:39.02" />
                    <SPLIT distance="900" swimtime="00:08:54.32" />
                    <SPLIT distance="925" swimtime="00:09:09.67" />
                    <SPLIT distance="950" swimtime="00:09:24.98" />
                    <SPLIT distance="975" swimtime="00:09:40.36" />
                    <SPLIT distance="1000" swimtime="00:09:55.71" />
                    <SPLIT distance="1025" swimtime="00:10:10.99" />
                    <SPLIT distance="1050" swimtime="00:10:26.30" />
                    <SPLIT distance="1075" swimtime="00:10:41.55" />
                    <SPLIT distance="1100" swimtime="00:10:56.93" />
                    <SPLIT distance="1125" swimtime="00:11:12.13" />
                    <SPLIT distance="1150" swimtime="00:11:27.60" />
                    <SPLIT distance="1175" swimtime="00:11:42.75" />
                    <SPLIT distance="1200" swimtime="00:11:58.06" />
                    <SPLIT distance="1225" swimtime="00:12:13.43" />
                    <SPLIT distance="1250" swimtime="00:12:28.58" />
                    <SPLIT distance="1275" swimtime="00:12:43.74" />
                    <SPLIT distance="1300" swimtime="00:12:58.99" />
                    <SPLIT distance="1325" swimtime="00:13:14.46" />
                    <SPLIT distance="1350" swimtime="00:13:29.77" />
                    <SPLIT distance="1375" swimtime="00:13:45.07" />
                    <SPLIT distance="1400" swimtime="00:14:00.38" />
                    <SPLIT distance="1425" swimtime="00:14:15.67" />
                    <SPLIT distance="1450" swimtime="00:14:30.49" />
                    <SPLIT distance="1475" swimtime="00:14:45.37" />
                    <SPLIT distance="1500" swimtime="00:14:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="11" lane="5" heat="1" heatid="10042" swimtime="00:07:44.53" reactiontime="+65" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="75" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:00:55.09" />
                    <SPLIT distance="125" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:23.85" />
                    <SPLIT distance="175" swimtime="00:01:38.39" />
                    <SPLIT distance="200" swimtime="00:01:52.91" />
                    <SPLIT distance="225" swimtime="00:02:07.31" />
                    <SPLIT distance="250" swimtime="00:02:21.67" />
                    <SPLIT distance="275" swimtime="00:02:36.16" />
                    <SPLIT distance="300" swimtime="00:02:50.79" />
                    <SPLIT distance="325" swimtime="00:03:05.46" />
                    <SPLIT distance="350" swimtime="00:03:20.11" />
                    <SPLIT distance="375" swimtime="00:03:34.81" />
                    <SPLIT distance="400" swimtime="00:03:49.37" />
                    <SPLIT distance="425" swimtime="00:04:03.92" />
                    <SPLIT distance="450" swimtime="00:04:18.65" />
                    <SPLIT distance="475" swimtime="00:04:33.35" />
                    <SPLIT distance="500" swimtime="00:04:48.05" />
                    <SPLIT distance="525" swimtime="00:05:02.81" />
                    <SPLIT distance="550" swimtime="00:05:17.51" />
                    <SPLIT distance="575" swimtime="00:05:32.30" />
                    <SPLIT distance="600" swimtime="00:05:47.05" />
                    <SPLIT distance="625" swimtime="00:06:01.87" />
                    <SPLIT distance="650" swimtime="00:06:16.59" />
                    <SPLIT distance="675" swimtime="00:06:31.43" />
                    <SPLIT distance="700" swimtime="00:06:46.25" />
                    <SPLIT distance="725" swimtime="00:07:01.04" />
                    <SPLIT distance="750" swimtime="00:07:15.95" />
                    <SPLIT distance="775" swimtime="00:07:30.61" />
                    <SPLIT distance="800" swimtime="00:07:44.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108847" lastname="GONZALEZ" firstname="Hugo" gender="M" birthdate="1999-02-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.22" eventid="46" heat="2" lane="3">
                  <MEETINFO date="2021-11-27" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.61" eventid="7" heat="4" lane="8">
                  <MEETINFO date="2021-07-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="12" lane="3" heat="2" heatid="20046" swimtime="00:01:52.02" reactiontime="+63" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                    <SPLIT distance="75" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:00:54.89" />
                    <SPLIT distance="125" swimtime="00:01:09.31" />
                    <SPLIT distance="150" swimtime="00:01:23.58" />
                    <SPLIT distance="175" swimtime="00:01:37.92" />
                    <SPLIT distance="200" swimtime="00:01:52.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="21" lane="8" heat="4" heatid="40007" swimtime="00:01:57.27" reactiontime="+64" points="817">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:25.25" />
                    <SPLIT distance="75" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:00:54.45" />
                    <SPLIT distance="125" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:28.12" />
                    <SPLIT distance="175" swimtime="00:01:43.14" />
                    <SPLIT distance="200" swimtime="00:01:57.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213230" lastname="DOMINGUEZ" firstname="Luis" gender="M" birthdate="2003-01-18">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.59" eventid="44" heat="3" lane="4">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:03:47.63" eventid="24" heat="2" lane="3">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="20" lane="4" heat="3" heatid="30044" swimtime="00:01:44.25" reactiontime="+68" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                    <SPLIT distance="75" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:00:49.72" />
                    <SPLIT distance="125" swimtime="00:01:03.10" />
                    <SPLIT distance="150" swimtime="00:01:16.76" />
                    <SPLIT distance="175" swimtime="00:01:30.54" />
                    <SPLIT distance="200" swimtime="00:01:44.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="16" lane="3" heat="2" heatid="20024" swimtime="00:03:43.18" reactiontime="+71" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.89" />
                    <SPLIT distance="75" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:00:52.48" />
                    <SPLIT distance="125" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:20.66" />
                    <SPLIT distance="175" swimtime="00:01:34.80" />
                    <SPLIT distance="200" swimtime="00:01:49.13" />
                    <SPLIT distance="225" swimtime="00:02:03.35" />
                    <SPLIT distance="250" swimtime="00:02:17.54" />
                    <SPLIT distance="275" swimtime="00:02:31.94" />
                    <SPLIT distance="300" swimtime="00:02:46.35" />
                    <SPLIT distance="325" swimtime="00:03:00.85" />
                    <SPLIT distance="350" swimtime="00:03:15.15" />
                    <SPLIT distance="375" swimtime="00:03:29.64" />
                    <SPLIT distance="400" swimtime="00:03:43.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124374" lastname="LOZANO" firstname="Alberto" gender="M" birthdate="1998-08-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:22.87" eventid="5" heat="7" lane="5">
                  <MEETINFO date="2021-11-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="44" lane="5" heat="7" heatid="70005" swimtime="00:00:23.43" reactiontime="+63" points="799">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108846" lastname="ZAMORANO SANZ" firstname="Africa" gender="F" birthdate="1998-01-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.79" eventid="2" heat="5" lane="8">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.37" eventid="45" heat="4" lane="7">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.50" eventid="22" heat="3" lane="2">
                  <MEETINFO date="2021-11-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="22" lane="8" heat="5" heatid="50002" swimtime="00:00:58.28" reactiontime="+55" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.79" />
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                    <SPLIT distance="75" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:00:58.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="11" lane="7" heat="4" heatid="40045" swimtime="00:02:04.85" reactiontime="+54" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="75" swimtime="00:00:45.28" />
                    <SPLIT distance="100" swimtime="00:01:01.34" />
                    <SPLIT distance="125" swimtime="00:01:17.48" />
                    <SPLIT distance="150" swimtime="00:01:33.66" />
                    <SPLIT distance="175" swimtime="00:01:49.49" />
                    <SPLIT distance="200" swimtime="00:02:04.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="14" lane="2" heat="3" heatid="30022" swimtime="00:00:59.99" reactiontime="+65" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="75" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:00:59.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="-1" lane="1" heat="1" heatid="10222" swimtime="00:01:00.00" status="DSQ" reactiontime="+66" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201566" lastname="OTERO FERNANDEZ" firstname="Paula" gender="F" birthdate="2004-03-30">
              <ENTRIES>
                <ENTRY entrytime="00:04:08.95" eventid="1" heat="2" lane="3">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="00:08:34.90" eventid="12" heat="2" lane="1">
                  <MEETINFO date="2022-04-09" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="20" lane="3" heat="2" heatid="20001" swimtime="00:04:14.08" reactiontime="+72" points="780">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="75" swimtime="00:00:44.04" />
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                    <SPLIT distance="125" swimtime="00:01:15.08" />
                    <SPLIT distance="150" swimtime="00:01:30.90" />
                    <SPLIT distance="175" swimtime="00:01:46.77" />
                    <SPLIT distance="200" swimtime="00:02:03.00" />
                    <SPLIT distance="225" swimtime="00:02:19.16" />
                    <SPLIT distance="250" swimtime="00:02:35.48" />
                    <SPLIT distance="275" swimtime="00:02:51.95" />
                    <SPLIT distance="300" swimtime="00:03:08.45" />
                    <SPLIT distance="325" swimtime="00:03:25.03" />
                    <SPLIT distance="350" swimtime="00:03:41.84" />
                    <SPLIT distance="375" swimtime="00:03:58.18" />
                    <SPLIT distance="400" swimtime="00:04:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="14" lane="1" heat="2" heatid="20012" swimtime="00:08:37.61" reactiontime="+73" points="794">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="75" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:01.66" />
                    <SPLIT distance="125" swimtime="00:01:17.66" />
                    <SPLIT distance="150" swimtime="00:01:33.58" />
                    <SPLIT distance="175" swimtime="00:01:49.49" />
                    <SPLIT distance="200" swimtime="00:02:05.40" />
                    <SPLIT distance="225" swimtime="00:02:21.15" />
                    <SPLIT distance="250" swimtime="00:02:37.01" />
                    <SPLIT distance="275" swimtime="00:02:52.77" />
                    <SPLIT distance="300" swimtime="00:03:08.77" />
                    <SPLIT distance="325" swimtime="00:03:24.76" />
                    <SPLIT distance="350" swimtime="00:03:41.00" />
                    <SPLIT distance="375" swimtime="00:03:57.14" />
                    <SPLIT distance="400" swimtime="00:04:13.53" />
                    <SPLIT distance="425" swimtime="00:04:29.60" />
                    <SPLIT distance="450" swimtime="00:04:46.01" />
                    <SPLIT distance="475" swimtime="00:05:02.34" />
                    <SPLIT distance="500" swimtime="00:05:18.80" />
                    <SPLIT distance="525" swimtime="00:05:35.34" />
                    <SPLIT distance="550" swimtime="00:05:52.00" />
                    <SPLIT distance="575" swimtime="00:06:08.47" />
                    <SPLIT distance="600" swimtime="00:06:25.25" />
                    <SPLIT distance="625" swimtime="00:06:41.95" />
                    <SPLIT distance="650" swimtime="00:06:58.71" />
                    <SPLIT distance="675" swimtime="00:07:15.32" />
                    <SPLIT distance="700" swimtime="00:07:32.12" />
                    <SPLIT distance="725" swimtime="00:07:48.75" />
                    <SPLIT distance="750" swimtime="00:08:05.52" />
                    <SPLIT distance="775" swimtime="00:08:21.91" />
                    <SPLIT distance="800" swimtime="00:08:37.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Spain">
              <RESULTS>
                <RESULT eventid="109" place="6" lane="2" heat="1" swimtime="00:03:07.19" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.86" />
                    <SPLIT distance="50" swimtime="00:00:22.70" />
                    <SPLIT distance="75" swimtime="00:00:34.83" />
                    <SPLIT distance="100" swimtime="00:00:46.90" />
                    <SPLIT distance="125" swimtime="00:00:57.27" />
                    <SPLIT distance="150" swimtime="00:01:09.13" />
                    <SPLIT distance="175" swimtime="00:01:21.37" />
                    <SPLIT distance="200" swimtime="00:01:33.53" />
                    <SPLIT distance="225" swimtime="00:01:43.63" />
                    <SPLIT distance="250" swimtime="00:01:55.21" />
                    <SPLIT distance="275" swimtime="00:02:07.38" />
                    <SPLIT distance="300" swimtime="00:02:19.97" />
                    <SPLIT distance="325" swimtime="00:02:30.19" />
                    <SPLIT distance="350" swimtime="00:02:42.11" />
                    <SPLIT distance="375" swimtime="00:02:54.57" />
                    <SPLIT distance="400" swimtime="00:03:07.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154217" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="213230" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="182683" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="154214" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="5" lane="6" heat="1" swimtime="00:03:07.75" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.74" />
                    <SPLIT distance="50" swimtime="00:00:22.53" />
                    <SPLIT distance="75" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:00:46.71" />
                    <SPLIT distance="125" swimtime="00:00:56.76" />
                    <SPLIT distance="150" swimtime="00:01:08.59" />
                    <SPLIT distance="175" swimtime="00:01:20.84" />
                    <SPLIT distance="200" swimtime="00:01:33.08" />
                    <SPLIT distance="225" swimtime="00:01:43.38" />
                    <SPLIT distance="250" swimtime="00:01:55.26" />
                    <SPLIT distance="275" swimtime="00:02:07.40" />
                    <SPLIT distance="300" swimtime="00:02:19.77" />
                    <SPLIT distance="325" swimtime="00:02:30.39" />
                    <SPLIT distance="350" swimtime="00:02:42.77" />
                    <SPLIT distance="375" swimtime="00:02:55.31" />
                    <SPLIT distance="400" swimtime="00:03:07.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154217" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="213230" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="182683" reactiontime="+21" />
                    <RELAYPOSITION number="4" athleteid="154214" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Spain">
              <RESULTS>
                <RESULT eventid="48" place="9" lane="1" heat="2" swimtime="00:03:26.48" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.28" />
                    <SPLIT distance="75" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:00:51.86" />
                    <SPLIT distance="125" swimtime="00:01:03.79" />
                    <SPLIT distance="150" swimtime="00:01:18.81" />
                    <SPLIT distance="175" swimtime="00:01:34.23" />
                    <SPLIT distance="200" swimtime="00:01:50.10" />
                    <SPLIT distance="225" swimtime="00:02:00.37" />
                    <SPLIT distance="250" swimtime="00:02:13.33" />
                    <SPLIT distance="275" swimtime="00:02:26.72" />
                    <SPLIT distance="300" swimtime="00:02:40.46" />
                    <SPLIT distance="325" swimtime="00:02:50.86" />
                    <SPLIT distance="350" swimtime="00:03:02.61" />
                    <SPLIT distance="375" swimtime="00:03:14.58" />
                    <SPLIT distance="400" swimtime="00:03:26.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="108847" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="154214" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="182683" reactiontime="+1" />
                    <RELAYPOSITION number="4" athleteid="154217" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Spain">
              <RESULTS>
                <RESULT eventid="132" place="6" lane="1" heat="1" swimtime="00:06:53.13" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.20" />
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                    <SPLIT distance="75" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:00:49.46" />
                    <SPLIT distance="125" swimtime="00:01:02.67" />
                    <SPLIT distance="150" swimtime="00:01:16.16" />
                    <SPLIT distance="175" swimtime="00:01:29.84" />
                    <SPLIT distance="200" swimtime="00:01:43.02" />
                    <SPLIT distance="225" swimtime="00:01:53.31" />
                    <SPLIT distance="250" swimtime="00:02:05.68" />
                    <SPLIT distance="275" swimtime="00:02:18.39" />
                    <SPLIT distance="300" swimtime="00:02:31.40" />
                    <SPLIT distance="325" swimtime="00:02:44.60" />
                    <SPLIT distance="350" swimtime="00:02:58.31" />
                    <SPLIT distance="375" swimtime="00:03:12.22" />
                    <SPLIT distance="400" swimtime="00:03:25.71" />
                    <SPLIT distance="425" swimtime="00:03:36.63" />
                    <SPLIT distance="450" swimtime="00:03:49.34" />
                    <SPLIT distance="475" swimtime="00:04:02.34" />
                    <SPLIT distance="500" swimtime="00:04:15.65" />
                    <SPLIT distance="525" swimtime="00:04:29.06" />
                    <SPLIT distance="550" swimtime="00:04:42.98" />
                    <SPLIT distance="575" swimtime="00:04:56.69" />
                    <SPLIT distance="600" swimtime="00:05:10.01" />
                    <SPLIT distance="625" swimtime="00:05:20.82" />
                    <SPLIT distance="650" swimtime="00:05:33.36" />
                    <SPLIT distance="675" swimtime="00:05:46.38" />
                    <SPLIT distance="700" swimtime="00:05:59.56" />
                    <SPLIT distance="725" swimtime="00:06:12.78" />
                    <SPLIT distance="750" swimtime="00:06:26.17" />
                    <SPLIT distance="775" swimtime="00:06:39.84" />
                    <SPLIT distance="800" swimtime="00:06:53.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213230" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="182683" reactiontime="+12" />
                    <RELAYPOSITION number="3" athleteid="108847" reactiontime="+16" />
                    <RELAYPOSITION number="4" athleteid="154217" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="7" lane="2" heat="1" swimtime="00:06:56.79" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:24.40" />
                    <SPLIT distance="75" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:00:50.96" />
                    <SPLIT distance="125" swimtime="00:01:04.32" />
                    <SPLIT distance="150" swimtime="00:01:17.98" />
                    <SPLIT distance="175" swimtime="00:01:31.71" />
                    <SPLIT distance="200" swimtime="00:01:45.16" />
                    <SPLIT distance="225" swimtime="00:01:55.76" />
                    <SPLIT distance="250" swimtime="00:02:08.05" />
                    <SPLIT distance="275" swimtime="00:02:20.87" />
                    <SPLIT distance="300" swimtime="00:02:34.01" />
                    <SPLIT distance="325" swimtime="00:02:47.48" />
                    <SPLIT distance="350" swimtime="00:03:01.33" />
                    <SPLIT distance="375" swimtime="00:03:15.14" />
                    <SPLIT distance="400" swimtime="00:03:28.67" />
                    <SPLIT distance="425" swimtime="00:03:39.32" />
                    <SPLIT distance="450" swimtime="00:03:52.39" />
                    <SPLIT distance="475" swimtime="00:04:05.44" />
                    <SPLIT distance="500" swimtime="00:04:18.55" />
                    <SPLIT distance="525" swimtime="00:04:31.97" />
                    <SPLIT distance="550" swimtime="00:04:45.39" />
                    <SPLIT distance="575" swimtime="00:04:59.08" />
                    <SPLIT distance="600" swimtime="00:05:12.24" />
                    <SPLIT distance="625" swimtime="00:05:23.23" />
                    <SPLIT distance="650" swimtime="00:05:36.08" />
                    <SPLIT distance="675" swimtime="00:05:49.18" />
                    <SPLIT distance="700" swimtime="00:06:02.52" />
                    <SPLIT distance="725" swimtime="00:06:15.95" />
                    <SPLIT distance="750" swimtime="00:06:29.46" />
                    <SPLIT distance="775" swimtime="00:06:43.09" />
                    <SPLIT distance="800" swimtime="00:06:56.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154217" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="182683" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="213230" reactiontime="+16" />
                    <RELAYPOSITION number="4" athleteid="108847" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Spain">
              <RESULTS>
                <RESULT eventid="126" place="6" lane="1" heat="1" swimtime="00:01:24.83" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.32" />
                    <SPLIT distance="50" swimtime="00:00:21.59" />
                    <SPLIT distance="75" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:00:42.67" />
                    <SPLIT distance="125" swimtime="00:00:52.74" />
                    <SPLIT distance="150" swimtime="00:01:03.71" />
                    <SPLIT distance="175" swimtime="00:01:13.60" />
                    <SPLIT distance="200" swimtime="00:01:24.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154214" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="213230" reactiontime="+11" />
                    <RELAYPOSITION number="3" athleteid="154217" reactiontime="+15" />
                    <RELAYPOSITION number="4" athleteid="182683" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="7" lane="8" heat="2" swimtime="00:01:26.29" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:21.78" />
                    <SPLIT distance="75" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:00:43.30" />
                    <SPLIT distance="125" swimtime="00:00:53.57" />
                    <SPLIT distance="150" swimtime="00:01:05.02" />
                    <SPLIT distance="175" swimtime="00:01:14.95" />
                    <SPLIT distance="200" swimtime="00:01:26.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154214" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="154217" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="182683" reactiontime="+17" />
                    <RELAYPOSITION number="4" athleteid="213230" reactiontime="-2" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Spain">
              <RESULTS>
                <RESULT eventid="35" place="-1" lane="7" heat="1" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Estonia" shortname="EST" code="EST" nation="EST" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="141785" lastname="LELLE" firstname="Armin Evert" gender="M" birthdate="1999-06-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.00" eventid="3" heat="5" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.20" eventid="46" heat="4" lane="2">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.52" eventid="19" heat="3" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="25" lane="2" heat="5" heatid="50003" swimtime="00:00:52.39" reactiontime="+63" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:25.26" />
                    <SPLIT distance="75" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:00:52.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="20" lane="2" heat="4" heatid="40046" swimtime="00:01:54.16" reactiontime="+64" points="792">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.83" />
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                    <SPLIT distance="75" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:00:55.48" />
                    <SPLIT distance="125" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:24.69" />
                    <SPLIT distance="175" swimtime="00:01:39.58" />
                    <SPLIT distance="200" swimtime="00:01:54.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="34" lane="7" heat="3" heatid="30019" swimtime="00:00:24.69" reactiontime="+65" points="728">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                    <SPLIT distance="50" swimtime="00:00:24.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="137206" lastname="ZAITSEV" firstname="Daniel" gender="M" birthdate="1997-12-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.50" eventid="39" heat="7" lane="8">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.08" eventid="14" heat="9" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.51" eventid="5" heat="10" lane="2">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.38" eventid="31" heat="9" lane="8">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="14" lane="8" heat="7" heatid="70039" swimtime="00:00:50.55" reactiontime="+68" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.56" />
                    <SPLIT distance="50" swimtime="00:00:23.41" />
                    <SPLIT distance="75" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:00:50.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="12" lane="1" heat="1" heatid="10239" swimtime="00:00:50.48" reactiontime="+65" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.32" />
                    <SPLIT distance="50" swimtime="00:00:22.99" />
                    <SPLIT distance="75" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:00:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="29" lane="1" heat="9" heatid="90014" swimtime="00:00:47.46" reactiontime="+67" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.53" />
                    <SPLIT distance="50" swimtime="00:00:22.58" />
                    <SPLIT distance="75" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:00:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="105" place="8" lane="8" heat="1" heatid="10105" swimtime="00:00:22.38" reactiontime="+64" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="12" lane="2" heat="10" heatid="100005" swimtime="00:00:22.41" reactiontime="+64" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.19" />
                    <SPLIT distance="50" swimtime="00:00:22.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="8" lane="7" heat="1" heatid="10205" swimtime="00:00:22.28" reactiontime="+60" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.07" />
                    <SPLIT distance="50" swimtime="00:00:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="405" place="8" lane="5" heat="1" heatid="10405" swimtime="00:00:22.15" reactiontime="+59" points="946">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.03" />
                    <SPLIT distance="50" swimtime="00:00:22.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="18" lane="8" heat="9" heatid="90031" swimtime="00:00:21.33" reactiontime="+64" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="331" place="19" lane="3" heat="1" heatid="10331" swimtime="00:00:21.34" reactiontime="+63" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:21.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108611" lastname="ZIRK" firstname="Kregor" gender="M" birthdate="1999-07-03">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.68" eventid="21" heat="3" lane="3">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.58" eventid="44" heat="5" lane="1">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="121" place="5" lane="7" heat="1" heatid="10121" swimtime="00:01:50.51" reactiontime="+63" points="939">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.21" />
                    <SPLIT distance="50" swimtime="00:00:24.72" />
                    <SPLIT distance="75" swimtime="00:00:38.70" />
                    <SPLIT distance="100" swimtime="00:00:52.75" />
                    <SPLIT distance="125" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:21.47" />
                    <SPLIT distance="175" swimtime="00:01:36.11" />
                    <SPLIT distance="200" swimtime="00:01:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="6" lane="3" heat="3" heatid="30021" swimtime="00:01:50.85" reactiontime="+63" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.26" />
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="75" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:00:53.17" />
                    <SPLIT distance="125" swimtime="00:01:07.47" />
                    <SPLIT distance="150" swimtime="00:01:22.00" />
                    <SPLIT distance="175" swimtime="00:01:36.48" />
                    <SPLIT distance="200" swimtime="00:01:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="11" lane="1" heat="5" heatid="50044" swimtime="00:01:43.16" reactiontime="+59" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.30" />
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="75" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:00:50.55" />
                    <SPLIT distance="125" swimtime="00:01:03.75" />
                    <SPLIT distance="150" swimtime="00:01:17.00" />
                    <SPLIT distance="175" swimtime="00:01:30.38" />
                    <SPLIT distance="200" swimtime="00:01:43.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100393" lastname="ROMANJUK" firstname="Maria" gender="F" birthdate="1996-08-15">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.93" eventid="15" heat="4" lane="8">
                  <MEETINFO date="2021-10-08" />
                </ENTRY>
                <ENTRY entrytime="00:02:25.95" eventid="28" heat="2" lane="6">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.32" eventid="6" heat="2" lane="7">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.30" eventid="40" heat="4" lane="7">
                  <MEETINFO date="2021-11-26" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.24" eventid="22" heat="2" lane="1">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="25" lane="8" heat="4" heatid="40015" swimtime="00:01:06.26" reactiontime="+68" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.35" />
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="75" swimtime="00:00:48.56" />
                    <SPLIT distance="100" swimtime="00:01:06.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="23" lane="6" heat="2" heatid="20028" swimtime="00:02:25.53" reactiontime="+69" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="75" swimtime="00:00:50.93" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="125" swimtime="00:01:28.28" />
                    <SPLIT distance="150" swimtime="00:01:47.20" />
                    <SPLIT distance="175" swimtime="00:02:06.47" />
                    <SPLIT distance="200" swimtime="00:02:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="31" lane="7" heat="2" heatid="20006" swimtime="00:02:14.15" reactiontime="+69" points="749">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="75" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                    <SPLIT distance="125" swimtime="00:01:22.88" />
                    <SPLIT distance="150" swimtime="00:01:42.19" />
                    <SPLIT distance="175" swimtime="00:01:59.02" />
                    <SPLIT distance="200" swimtime="00:02:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="-1" lane="7" heat="4" heatid="40040" swimtime="00:00:30.99" status="DSQ" reactiontime="+67" />
                <RESULT eventid="22" place="19" lane="1" heat="2" heatid="20022" swimtime="00:01:01.32" reactiontime="+65" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                    <SPLIT distance="75" swimtime="00:00:46.10" />
                    <SPLIT distance="100" swimtime="00:01:01.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Fiji" shortname="FIJ" code="FIJ" nation="FIJ" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="180567" lastname="MCCAIG" firstname="Hansel" gender="M" birthdate="2003-07-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.40" eventid="14" heat="5" lane="8">
                  <MEETINFO date="2022-07-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.29" eventid="31" heat="5" lane="2">
                  <MEETINFO date="2022-08-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="49" lane="8" heat="5" heatid="50014" swimtime="00:00:49.73" reactiontime="+58" points="733">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.10" />
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="75" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:00:49.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="49" lane="2" heat="5" heatid="50031" swimtime="00:00:22.61" reactiontime="+58" points="708">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.86" />
                    <SPLIT distance="50" swimtime="00:00:22.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123169" lastname="RABUA" firstname="Epeli Herbert Jordan" gender="M" birthdate="1998-10-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.60" eventid="41" heat="3" lane="1">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.01" eventid="5" heat="3" lane="3">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="49" lane="1" heat="3" heatid="30041" swimtime="00:00:28.84" reactiontime="+63" points="647">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="54" lane="3" heat="3" heatid="30005" swimtime="00:00:25.60" reactiontime="+66" points="613">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.79" />
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201784" lastname="MUDUNASOKO" firstname="Kelera" gender="F" birthdate="2007-07-20">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.94" eventid="15" heat="2" lane="8">
                  <MEETINFO date="2022-04-09" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.14" eventid="40" heat="3" lane="2">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="44" lane="8" heat="2" heatid="20015" swimtime="00:01:13.86" reactiontime="+70" points="601">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.00" />
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="75" swimtime="00:00:53.98" />
                    <SPLIT distance="100" swimtime="00:01:13.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="34" lane="2" heat="3" heatid="30040" swimtime="00:00:34.05" reactiontime="+67" points="590">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149586" lastname="ROVA" firstname="Rosemarie" gender="F" birthdate="2002-09-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.90" eventid="4" heat="2" lane="5">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.08" eventid="30" heat="3" lane="3">
                  <MEETINFO date="2022-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="-1" lane="5" heat="2" heatid="20004" swimtime="NT" status="DNS" />
                <RESULT eventid="30" place="-1" lane="3" heat="3" heatid="30030" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Finland" shortname="FIN" code="FIN" nation="FIN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198386" lastname="KOKKO" firstname="Olli" gender="M" birthdate="1994-04-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.04" eventid="16" heat="5" lane="5">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.35" eventid="41" heat="9" lane="7">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="-1" lane="5" heat="5" heatid="50016" swimtime="00:00:58.15" status="DSQ" reactiontime="+64" />
                <RESULT eventid="41" place="16" lane="7" heat="9" heatid="90041" swimtime="00:00:26.51" reactiontime="+65" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.00" />
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="11" lane="8" heat="1" heatid="10241" swimtime="00:00:26.25" reactiontime="+64" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="341" place="16" lane="5" heat="1" heatid="10341" swimtime="00:00:26.24" reactiontime="+59" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191727" lastname="BRÄNNKÄRR" firstname="Ronny" gender="M" birthdate="2002-07-11">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.90" eventid="44" heat="3" lane="6">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:01:56.59" eventid="7" heat="5" lane="1">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.68" eventid="23" heat="5" lane="7">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="26" lane="6" heat="3" heatid="30044" swimtime="00:01:45.42" reactiontime="+67" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                    <SPLIT distance="75" swimtime="00:00:37.85" />
                    <SPLIT distance="100" swimtime="00:00:51.54" />
                    <SPLIT distance="125" swimtime="00:01:04.90" />
                    <SPLIT distance="150" swimtime="00:01:18.36" />
                    <SPLIT distance="175" swimtime="00:01:31.93" />
                    <SPLIT distance="200" swimtime="00:01:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="19" lane="1" heat="5" heatid="50007" swimtime="00:01:55.33" reactiontime="+65" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.78" />
                    <SPLIT distance="50" swimtime="00:00:24.12" />
                    <SPLIT distance="75" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:00:52.95" />
                    <SPLIT distance="125" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:26.93" />
                    <SPLIT distance="175" swimtime="00:01:41.49" />
                    <SPLIT distance="200" swimtime="00:01:55.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="17" lane="7" heat="5" heatid="50023" swimtime="00:00:52.81" reactiontime="+68" points="812">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.59" />
                    <SPLIT distance="75" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:00:52.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="323" place="18" lane="5" heat="1" heatid="10323" swimtime="00:00:52.28" reactiontime="+65" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.56" />
                    <SPLIT distance="50" swimtime="00:00:23.45" />
                    <SPLIT distance="75" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:00:52.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100849" lastname="KIVIRINTA" firstname="Veera" gender="F" birthdate="1995-04-06">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.44" eventid="15" heat="5" lane="1">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.85" eventid="40" heat="6" lane="6">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="30" lane="1" heat="5" heatid="50015" swimtime="00:01:06.59" reactiontime="+73" points="821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="75" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="8" lane="8" heat="1" heatid="10140" swimtime="00:00:29.84" reactiontime="+74" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="8" lane="6" heat="6" heatid="60040" swimtime="00:00:29.72" reactiontime="+75" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="8" lane="6" heat="1" heatid="10240" swimtime="00:00:29.80" reactiontime="+75" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157490" lastname="HULKKO" firstname="Ida" gender="F" birthdate="1998-12-12">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.98" eventid="15" heat="7" lane="2">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.62" eventid="40" heat="5" lane="3">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="14" lane="2" heat="7" heatid="70015" swimtime="00:01:05.25" reactiontime="+67" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.79" />
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="75" swimtime="00:00:47.56" />
                    <SPLIT distance="100" swimtime="00:01:05.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="9" lane="1" heat="1" heatid="10215" swimtime="00:01:04.85" reactiontime="+66" points="889">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="75" swimtime="00:00:47.21" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="12" lane="3" heat="5" heatid="50040" swimtime="00:00:29.89" reactiontime="+64" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="10" lane="7" heat="1" heatid="10240" swimtime="00:00:29.94" reactiontime="+65" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166204" lastname="LAHTINEN" firstname="Laura" gender="F" birthdate="2003-06-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.13" eventid="38" heat="3" lane="2">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.78" eventid="28" heat="2" lane="5">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.61" eventid="20" heat="3" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.97" eventid="43" heat="4" lane="1">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.76" eventid="6" heat="2" lane="4">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="16" lane="2" heat="3" heatid="30038" swimtime="00:00:57.85" reactiontime="+68" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                    <SPLIT distance="75" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:00:57.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="16" lane="8" heat="1" heatid="10238" swimtime="00:00:58.09" reactiontime="+68" points="829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                    <SPLIT distance="75" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:00:58.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="338" place="16" lane="5" heat="1" heatid="10338" swimtime="00:00:56.88" reactiontime="+68" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                    <SPLIT distance="75" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:00:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="27" lane="5" heat="2" heatid="20028" swimtime="00:02:28.80" reactiontime="+70" points="739">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.96" />
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="75" swimtime="00:00:50.55" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="125" swimtime="00:01:28.31" />
                    <SPLIT distance="150" swimtime="00:01:48.03" />
                    <SPLIT distance="175" swimtime="00:02:08.34" />
                    <SPLIT distance="200" swimtime="00:02:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="120" place="8" lane="6" heat="1" heatid="10120" swimtime="00:02:06.48" reactiontime="+68" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.76" />
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="75" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:00:59.76" />
                    <SPLIT distance="125" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:32.68" />
                    <SPLIT distance="175" swimtime="00:01:49.51" />
                    <SPLIT distance="200" swimtime="00:02:06.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="4" lane="3" heat="3" heatid="30020" swimtime="00:02:05.13" reactiontime="+70" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                    <SPLIT distance="75" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:00:59.64" />
                    <SPLIT distance="125" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:32.04" />
                    <SPLIT distance="175" swimtime="00:01:48.50" />
                    <SPLIT distance="200" swimtime="00:02:05.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="-1" lane="1" heat="4" heatid="40043" swimtime="NT" status="DNS" />
                <RESULT eventid="6" place="21" lane="4" heat="2" heatid="20006" swimtime="00:02:10.66" reactiontime="+69" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:01:00.52" />
                    <SPLIT distance="125" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:01:38.46" />
                    <SPLIT distance="175" swimtime="00:01:55.09" />
                    <SPLIT distance="200" swimtime="00:02:10.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="France" shortname="FRA" code="FRA" nation="FRA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="181969" lastname="TOMAC" firstname="Mewen" gender="M" birthdate="2001-09-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.06" eventid="3" heat="5" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.14" eventid="46" heat="4" lane="3">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.27" eventid="19" heat="5" lane="6">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="7" lane="8" heat="1" heatid="10103" swimtime="00:00:49.94" reactiontime="+57" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.10" />
                    <SPLIT distance="75" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:00:49.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="2" lane="3" heat="5" heatid="50003" swimtime="00:00:49.99" reactiontime="+59" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:24.01" />
                    <SPLIT distance="75" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:00:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="7" lane="4" heat="1" heatid="10203" swimtime="00:00:50.01" reactiontime="+59" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:23.89" />
                    <SPLIT distance="75" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="146" place="6" lane="5" heat="1" heatid="10146" swimtime="00:01:49.93" reactiontime="+63" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:25.44" />
                    <SPLIT distance="75" swimtime="00:00:39.21" />
                    <SPLIT distance="100" swimtime="00:00:53.22" />
                    <SPLIT distance="125" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:21.80" />
                    <SPLIT distance="175" swimtime="00:01:35.97" />
                    <SPLIT distance="200" swimtime="00:01:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="2" lane="3" heat="4" heatid="40046" swimtime="00:01:49.61" reactiontime="+59" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                    <SPLIT distance="75" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:00:53.19" />
                    <SPLIT distance="125" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:21.42" />
                    <SPLIT distance="175" swimtime="00:01:35.67" />
                    <SPLIT distance="200" swimtime="00:01:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="20" lane="6" heat="5" heatid="50019" swimtime="00:00:23.58" reactiontime="+57" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:23.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191730" lastname="NDOYE-BROUARD" firstname="Yohann" gender="M" birthdate="2000-11-29">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.54" eventid="3" heat="6" lane="6">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.53" eventid="46" heat="4" lane="6">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="8" lane="2" heat="1" heatid="10103" swimtime="00:00:50.01" reactiontime="+60" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:24.17" />
                    <SPLIT distance="75" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="8" lane="6" heat="6" heatid="60003" swimtime="00:00:50.21" reactiontime="+56" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:24.04" />
                    <SPLIT distance="75" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:00:50.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="5" lane="6" heat="1" heatid="10203" swimtime="00:00:49.78" reactiontime="+59" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:24.28" />
                    <SPLIT distance="75" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:00:49.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="146" place="4" lane="2" heat="1" heatid="10146" swimtime="00:01:49.23" reactiontime="+61" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:25.12" />
                    <SPLIT distance="75" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:00:52.31" />
                    <SPLIT distance="125" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:20.13" />
                    <SPLIT distance="175" swimtime="00:01:34.56" />
                    <SPLIT distance="200" swimtime="00:01:49.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="5" lane="6" heat="4" heatid="40046" swimtime="00:01:50.12" reactiontime="+60" points="882">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.95" />
                    <SPLIT distance="50" swimtime="00:00:25.44" />
                    <SPLIT distance="75" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:00:53.01" />
                    <SPLIT distance="125" swimtime="00:01:07.18" />
                    <SPLIT distance="150" swimtime="00:01:21.82" />
                    <SPLIT distance="175" swimtime="00:01:36.30" />
                    <SPLIT distance="200" swimtime="00:01:50.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197601" lastname="VIQUERAT" firstname="Antoine" gender="M" birthdate="1998-10-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.53" eventid="16" heat="7" lane="7">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.86" eventid="29" heat="3" lane="6">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="5" lane="8" heat="1" heatid="10116" swimtime="00:00:56.98" reactiontime="+69" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                    <SPLIT distance="75" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:00:56.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="7" lane="7" heat="7" heatid="70016" swimtime="00:00:57.18" reactiontime="+67" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="75" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:00:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="8" lane="6" heat="2" heatid="20216" swimtime="00:00:57.07" reactiontime="+69" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:00:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="129" place="6" lane="2" heat="1" heatid="10129" swimtime="00:02:03.33" reactiontime="+66" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                    <SPLIT distance="75" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:00:59.53" />
                    <SPLIT distance="125" swimtime="00:01:15.54" />
                    <SPLIT distance="150" swimtime="00:01:31.45" />
                    <SPLIT distance="175" swimtime="00:01:47.39" />
                    <SPLIT distance="200" swimtime="00:02:03.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="5" lane="6" heat="3" heatid="30029" swimtime="00:02:03.93" reactiontime="+74" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                    <SPLIT distance="75" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="125" swimtime="00:01:15.81" />
                    <SPLIT distance="150" swimtime="00:01:31.79" />
                    <SPLIT distance="175" swimtime="00:01:47.67" />
                    <SPLIT distance="200" swimtime="00:02:03.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201991" lastname="AIT KACI" firstname="Carl" gender="M" birthdate="2001-06-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.58" eventid="16" heat="6" lane="1">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.47" eventid="29" heat="3" lane="2">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.70" eventid="41" heat="9" lane="8">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="12" lane="1" heat="6" heatid="60016" swimtime="00:00:57.68" reactiontime="+67" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.03" />
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                    <SPLIT distance="75" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:00:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="16" lane="7" heat="1" heatid="10216" swimtime="00:00:58.12" reactiontime="+69" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                    <SPLIT distance="75" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:00:58.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="-1" lane="2" heat="3" heatid="30029" swimtime="00:02:06.39" status="DSQ" reactiontime="+75" />
                <RESULT eventid="41" place="11" lane="8" heat="9" heatid="90041" swimtime="00:00:26.37" reactiontime="+62" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:26.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="14" lane="7" heat="1" heatid="10241" swimtime="00:00:26.41" reactiontime="+62" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149769" lastname="GROUSSET" firstname="Maxime" gender="M" birthdate="1999-04-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.61" eventid="14" heat="9" lane="4">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.09" eventid="44" heat="5" lane="3">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.03" eventid="31" heat="11" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:51.49" eventid="23" heat="4" lane="5">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="2" lane="5" heat="1" heatid="10114" swimtime="00:00:45.41" reactiontime="+62" points="962">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.67" />
                    <SPLIT distance="75" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:00:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="2" lane="4" heat="9" heatid="90014" swimtime="00:00:45.77" reactiontime="+63" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.38" />
                    <SPLIT distance="50" swimtime="00:00:21.85" />
                    <SPLIT distance="75" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:00:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="2" lane="4" heat="1" heatid="10214" swimtime="00:00:45.58" reactiontime="+64" points="952">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.51" />
                    <SPLIT distance="50" swimtime="00:00:22.12" />
                    <SPLIT distance="75" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:00:45.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="144" place="6" lane="3" heat="1" heatid="10144" swimtime="00:01:41.56" reactiontime="+61" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.99" />
                    <SPLIT distance="50" swimtime="00:00:23.54" />
                    <SPLIT distance="75" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:00:49.16" />
                    <SPLIT distance="125" swimtime="00:01:02.21" />
                    <SPLIT distance="150" swimtime="00:01:15.39" />
                    <SPLIT distance="175" swimtime="00:01:28.63" />
                    <SPLIT distance="200" swimtime="00:01:41.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="3" lane="3" heat="5" heatid="50044" swimtime="00:01:41.79" reactiontime="+63" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.85" />
                    <SPLIT distance="50" swimtime="00:00:23.27" />
                    <SPLIT distance="75" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:00:48.94" />
                    <SPLIT distance="125" swimtime="00:01:02.15" />
                    <SPLIT distance="150" swimtime="00:01:15.32" />
                    <SPLIT distance="175" swimtime="00:01:28.62" />
                    <SPLIT distance="200" swimtime="00:01:41.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="131" place="5" lane="8" heat="1" heatid="10131" swimtime="00:00:20.90" reactiontime="+63" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.07" />
                    <SPLIT distance="50" swimtime="00:00:20.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="10" lane="3" heat="11" heatid="110031" swimtime="00:00:21.13" reactiontime="+63" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.28" />
                    <SPLIT distance="50" swimtime="00:00:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="8" lane="2" heat="1" heatid="10231" swimtime="00:00:20.97" reactiontime="+67" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:20.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="1" lane="5" heat="4" heatid="40023" swimtime="00:00:51.94" reactiontime="+62" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:23.91" />
                    <SPLIT distance="75" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:00:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="-1" lane="4" heat="2" heatid="20223" swimtime="00:00:51.09" status="DSQ" reactiontime="+63" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100735" lastname="JOLY" firstname="Damien" gender="M" birthdate="1992-06-04">
              <ENTRIES>
                <ENTRY entrytime="00:14:25.62" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="2" lane="3" heat="5" heatid="30110" swimtime="00:14:19.62" reactiontime="+70" points="956">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                    <SPLIT distance="75" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:00:55.79" />
                    <SPLIT distance="125" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:24.49" />
                    <SPLIT distance="175" swimtime="00:01:38.93" />
                    <SPLIT distance="200" swimtime="00:01:53.45" />
                    <SPLIT distance="225" swimtime="00:02:07.91" />
                    <SPLIT distance="250" swimtime="00:02:22.37" />
                    <SPLIT distance="275" swimtime="00:02:36.80" />
                    <SPLIT distance="300" swimtime="00:02:51.27" />
                    <SPLIT distance="325" swimtime="00:03:05.67" />
                    <SPLIT distance="350" swimtime="00:03:20.13" />
                    <SPLIT distance="375" swimtime="00:03:34.47" />
                    <SPLIT distance="400" swimtime="00:03:48.92" />
                    <SPLIT distance="425" swimtime="00:04:03.33" />
                    <SPLIT distance="450" swimtime="00:04:17.74" />
                    <SPLIT distance="475" swimtime="00:04:32.25" />
                    <SPLIT distance="500" swimtime="00:04:46.60" />
                    <SPLIT distance="525" swimtime="00:05:00.98" />
                    <SPLIT distance="550" swimtime="00:05:15.32" />
                    <SPLIT distance="575" swimtime="00:05:29.66" />
                    <SPLIT distance="600" swimtime="00:05:43.89" />
                    <SPLIT distance="625" swimtime="00:05:58.36" />
                    <SPLIT distance="650" swimtime="00:06:12.66" />
                    <SPLIT distance="675" swimtime="00:06:26.96" />
                    <SPLIT distance="700" swimtime="00:06:41.33" />
                    <SPLIT distance="725" swimtime="00:06:55.66" />
                    <SPLIT distance="750" swimtime="00:07:10.13" />
                    <SPLIT distance="775" swimtime="00:07:24.48" />
                    <SPLIT distance="800" swimtime="00:07:38.82" />
                    <SPLIT distance="825" swimtime="00:07:53.19" />
                    <SPLIT distance="850" swimtime="00:08:07.50" />
                    <SPLIT distance="875" swimtime="00:08:21.73" />
                    <SPLIT distance="900" swimtime="00:08:36.05" />
                    <SPLIT distance="925" swimtime="00:08:50.28" />
                    <SPLIT distance="950" swimtime="00:09:04.62" />
                    <SPLIT distance="975" swimtime="00:09:18.96" />
                    <SPLIT distance="1000" swimtime="00:09:33.35" />
                    <SPLIT distance="1025" swimtime="00:09:47.56" />
                    <SPLIT distance="1050" swimtime="00:10:01.89" />
                    <SPLIT distance="1075" swimtime="00:10:16.22" />
                    <SPLIT distance="1100" swimtime="00:10:30.62" />
                    <SPLIT distance="1125" swimtime="00:10:44.83" />
                    <SPLIT distance="1150" swimtime="00:10:59.22" />
                    <SPLIT distance="1175" swimtime="00:11:13.58" />
                    <SPLIT distance="1200" swimtime="00:11:28.03" />
                    <SPLIT distance="1225" swimtime="00:11:42.33" />
                    <SPLIT distance="1250" swimtime="00:11:56.77" />
                    <SPLIT distance="1275" swimtime="00:12:11.18" />
                    <SPLIT distance="1300" swimtime="00:12:25.53" />
                    <SPLIT distance="1325" swimtime="00:12:40.00" />
                    <SPLIT distance="1350" swimtime="00:12:54.53" />
                    <SPLIT distance="1375" swimtime="00:13:09.09" />
                    <SPLIT distance="1400" swimtime="00:13:23.48" />
                    <SPLIT distance="1425" swimtime="00:13:37.83" />
                    <SPLIT distance="1450" swimtime="00:13:52.09" />
                    <SPLIT distance="1475" swimtime="00:14:06.17" />
                    <SPLIT distance="1500" swimtime="00:14:19.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144435" lastname="FONTAINE" firstname="Logan" gender="M" birthdate="1999-03-25">
              <ENTRIES>
                <ENTRY entrytime="00:14:36.82" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.00" eventid="24" heat="5" lane="7">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:07:35.47" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="5" lane="8" heat="5" heatid="30110" swimtime="00:14:27.90" reactiontime="+77" points="929">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.64" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="75" swimtime="00:00:41.01" />
                    <SPLIT distance="100" swimtime="00:00:55.29" />
                    <SPLIT distance="125" swimtime="00:01:09.70" />
                    <SPLIT distance="150" swimtime="00:01:24.11" />
                    <SPLIT distance="175" swimtime="00:01:38.58" />
                    <SPLIT distance="200" swimtime="00:01:53.29" />
                    <SPLIT distance="225" swimtime="00:02:07.81" />
                    <SPLIT distance="250" swimtime="00:02:22.36" />
                    <SPLIT distance="275" swimtime="00:02:36.87" />
                    <SPLIT distance="300" swimtime="00:02:51.36" />
                    <SPLIT distance="325" swimtime="00:03:05.89" />
                    <SPLIT distance="350" swimtime="00:03:20.46" />
                    <SPLIT distance="375" swimtime="00:03:34.95" />
                    <SPLIT distance="400" swimtime="00:03:49.54" />
                    <SPLIT distance="425" swimtime="00:04:04.21" />
                    <SPLIT distance="450" swimtime="00:04:18.68" />
                    <SPLIT distance="475" swimtime="00:04:33.18" />
                    <SPLIT distance="500" swimtime="00:04:47.85" />
                    <SPLIT distance="525" swimtime="00:05:02.52" />
                    <SPLIT distance="550" swimtime="00:05:16.97" />
                    <SPLIT distance="575" swimtime="00:05:31.42" />
                    <SPLIT distance="600" swimtime="00:05:45.95" />
                    <SPLIT distance="625" swimtime="00:06:00.54" />
                    <SPLIT distance="650" swimtime="00:06:15.06" />
                    <SPLIT distance="675" swimtime="00:06:29.55" />
                    <SPLIT distance="700" swimtime="00:06:44.08" />
                    <SPLIT distance="725" swimtime="00:06:58.53" />
                    <SPLIT distance="750" swimtime="00:07:13.09" />
                    <SPLIT distance="775" swimtime="00:07:27.70" />
                    <SPLIT distance="800" swimtime="00:07:42.26" />
                    <SPLIT distance="825" swimtime="00:07:56.90" />
                    <SPLIT distance="850" swimtime="00:08:11.38" />
                    <SPLIT distance="875" swimtime="00:08:25.98" />
                    <SPLIT distance="900" swimtime="00:08:40.69" />
                    <SPLIT distance="925" swimtime="00:08:55.30" />
                    <SPLIT distance="950" swimtime="00:09:09.86" />
                    <SPLIT distance="975" swimtime="00:09:24.41" />
                    <SPLIT distance="1000" swimtime="00:09:38.94" />
                    <SPLIT distance="1025" swimtime="00:09:53.45" />
                    <SPLIT distance="1050" swimtime="00:10:07.88" />
                    <SPLIT distance="1075" swimtime="00:10:22.45" />
                    <SPLIT distance="1100" swimtime="00:10:37.01" />
                    <SPLIT distance="1125" swimtime="00:10:51.49" />
                    <SPLIT distance="1150" swimtime="00:11:06.09" />
                    <SPLIT distance="1175" swimtime="00:11:20.73" />
                    <SPLIT distance="1200" swimtime="00:11:35.29" />
                    <SPLIT distance="1225" swimtime="00:11:49.81" />
                    <SPLIT distance="1250" swimtime="00:12:04.31" />
                    <SPLIT distance="1275" swimtime="00:12:18.92" />
                    <SPLIT distance="1300" swimtime="00:12:33.50" />
                    <SPLIT distance="1325" swimtime="00:12:48.23" />
                    <SPLIT distance="1350" swimtime="00:13:02.66" />
                    <SPLIT distance="1375" swimtime="00:13:17.29" />
                    <SPLIT distance="1400" swimtime="00:13:31.82" />
                    <SPLIT distance="1425" swimtime="00:13:46.00" />
                    <SPLIT distance="1450" swimtime="00:14:00.28" />
                    <SPLIT distance="1475" swimtime="00:14:14.32" />
                    <SPLIT distance="1500" swimtime="00:14:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="11" lane="7" heat="5" heatid="50024" swimtime="00:03:39.84" reactiontime="+74" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                    <SPLIT distance="50" swimtime="00:00:25.79" />
                    <SPLIT distance="75" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:00:53.54" />
                    <SPLIT distance="125" swimtime="00:01:07.37" />
                    <SPLIT distance="150" swimtime="00:01:21.34" />
                    <SPLIT distance="175" swimtime="00:01:35.23" />
                    <SPLIT distance="200" swimtime="00:01:49.34" />
                    <SPLIT distance="225" swimtime="00:02:03.17" />
                    <SPLIT distance="250" swimtime="00:02:17.26" />
                    <SPLIT distance="275" swimtime="00:02:31.04" />
                    <SPLIT distance="300" swimtime="00:02:45.06" />
                    <SPLIT distance="325" swimtime="00:02:58.85" />
                    <SPLIT distance="350" swimtime="00:03:12.81" />
                    <SPLIT distance="375" swimtime="00:03:26.43" />
                    <SPLIT distance="400" swimtime="00:03:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="3" lane="3" heat="5" heatid="30142" swimtime="00:07:33.12" reactiontime="+77" points="937">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:26.22" />
                    <SPLIT distance="75" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:00:54.18" />
                    <SPLIT distance="125" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:22.62" />
                    <SPLIT distance="175" swimtime="00:01:36.90" />
                    <SPLIT distance="200" swimtime="00:01:51.25" />
                    <SPLIT distance="225" swimtime="00:02:05.45" />
                    <SPLIT distance="250" swimtime="00:02:19.76" />
                    <SPLIT distance="275" swimtime="00:02:34.00" />
                    <SPLIT distance="300" swimtime="00:02:48.22" />
                    <SPLIT distance="325" swimtime="00:03:02.59" />
                    <SPLIT distance="350" swimtime="00:03:17.03" />
                    <SPLIT distance="375" swimtime="00:03:31.37" />
                    <SPLIT distance="400" swimtime="00:03:45.94" />
                    <SPLIT distance="425" swimtime="00:04:00.06" />
                    <SPLIT distance="450" swimtime="00:04:14.42" />
                    <SPLIT distance="475" swimtime="00:04:28.70" />
                    <SPLIT distance="500" swimtime="00:04:43.18" />
                    <SPLIT distance="525" swimtime="00:04:57.46" />
                    <SPLIT distance="550" swimtime="00:05:11.85" />
                    <SPLIT distance="575" swimtime="00:05:26.18" />
                    <SPLIT distance="600" swimtime="00:05:40.66" />
                    <SPLIT distance="625" swimtime="00:05:54.81" />
                    <SPLIT distance="650" swimtime="00:06:09.19" />
                    <SPLIT distance="675" swimtime="00:06:23.24" />
                    <SPLIT distance="700" swimtime="00:06:37.50" />
                    <SPLIT distance="725" swimtime="00:06:51.54" />
                    <SPLIT distance="750" swimtime="00:07:05.69" />
                    <SPLIT distance="775" swimtime="00:07:19.57" />
                    <SPLIT distance="800" swimtime="00:07:33.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201992" lastname="FUCHS" firstname="Roman" gender="M" birthdate="1998-01-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:43.16" eventid="44" heat="6" lane="7">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.85" eventid="24" heat="4" lane="1">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="12" lane="7" heat="6" heatid="60044" swimtime="00:01:43.17" reactiontime="+63" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:23.98" />
                    <SPLIT distance="75" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:00:50.00" />
                    <SPLIT distance="125" swimtime="00:01:03.28" />
                    <SPLIT distance="150" swimtime="00:01:16.65" />
                    <SPLIT distance="175" swimtime="00:01:30.01" />
                    <SPLIT distance="200" swimtime="00:01:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="-1" lane="1" heat="4" heatid="40024" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197605" lastname="MATTENET" firstname="Emilien" gender="M" birthdate="2000-11-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.30" eventid="7" heat="3" lane="7">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:04:08.16" eventid="37" heat="3" lane="1">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="24" lane="7" heat="3" heatid="30007" swimtime="00:01:57.91" reactiontime="+75" points="803">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.81" />
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                    <SPLIT distance="75" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:00:55.78" />
                    <SPLIT distance="125" swimtime="00:01:12.96" />
                    <SPLIT distance="150" swimtime="00:01:30.31" />
                    <SPLIT distance="175" swimtime="00:01:44.93" />
                    <SPLIT distance="200" swimtime="00:01:57.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="10" lane="1" heat="3" heatid="30037" swimtime="00:04:08.06" reactiontime="+71" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                    <SPLIT distance="75" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:00:57.45" />
                    <SPLIT distance="125" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:29.18" />
                    <SPLIT distance="175" swimtime="00:01:44.82" />
                    <SPLIT distance="200" swimtime="00:01:59.96" />
                    <SPLIT distance="225" swimtime="00:02:17.71" />
                    <SPLIT distance="250" swimtime="00:02:35.56" />
                    <SPLIT distance="275" swimtime="00:02:53.19" />
                    <SPLIT distance="300" swimtime="00:03:11.07" />
                    <SPLIT distance="325" swimtime="00:03:26.01" />
                    <SPLIT distance="350" swimtime="00:03:40.17" />
                    <SPLIT distance="375" swimtime="00:03:54.48" />
                    <SPLIT distance="400" swimtime="00:04:08.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101299" lastname="MANAUDOU" firstname="Florent" gender="M" birthdate="1990-11-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:22.68" eventid="5" heat="8" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.05" eventid="31" heat="10" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="16" lane="7" heat="8" heatid="80005" swimtime="00:00:22.53" reactiontime="+63" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.10" />
                    <SPLIT distance="50" swimtime="00:00:22.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="12" lane="8" heat="1" heatid="10205" swimtime="00:00:22.37" reactiontime="+64" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.00" />
                    <SPLIT distance="50" swimtime="00:00:22.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="305" place="16" lane="4" heat="1" heatid="10305" swimtime="00:00:22.31" reactiontime="+64" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.99" />
                    <SPLIT distance="50" swimtime="00:00:22.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="131" place="6" lane="1" heat="1" heatid="10131" swimtime="00:00:20.91" reactiontime="+60" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.90" />
                    <SPLIT distance="50" swimtime="00:00:20.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="4" lane="3" heat="10" heatid="100031" swimtime="00:00:20.94" reactiontime="+65" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.93" />
                    <SPLIT distance="50" swimtime="00:00:20.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="7" lane="5" heat="1" heatid="10231" swimtime="00:00:20.95" reactiontime="+65" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.04" />
                    <SPLIT distance="50" swimtime="00:00:20.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110511" lastname="MAHIEU" firstname="Pauline" gender="F" birthdate="1999-03-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.30" eventid="2" heat="4" lane="2">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.26" eventid="45" heat="5" lane="6">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="8" lane="2" heat="4" heatid="40002" swimtime="00:00:56.88" reactiontime="+60" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                    <SPLIT distance="75" swimtime="00:00:42.21" />
                    <SPLIT distance="100" swimtime="00:00:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="13" lane="6" heat="1" heatid="10202" swimtime="00:00:57.43" reactiontime="+58" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="75" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:00:57.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="7" lane="2" heat="1" heatid="10145" swimtime="00:02:03.21" reactiontime="+63" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="75" swimtime="00:00:44.49" />
                    <SPLIT distance="100" swimtime="00:01:00.32" />
                    <SPLIT distance="125" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:32.10" />
                    <SPLIT distance="175" swimtime="00:01:47.94" />
                    <SPLIT distance="200" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="5" lane="6" heat="5" heatid="50045" swimtime="00:02:02.96" reactiontime="+61" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                    <SPLIT distance="75" swimtime="00:00:44.77" />
                    <SPLIT distance="100" swimtime="00:01:00.20" />
                    <SPLIT distance="125" swimtime="00:01:15.77" />
                    <SPLIT distance="150" swimtime="00:01:31.75" />
                    <SPLIT distance="175" swimtime="00:01:47.65" />
                    <SPLIT distance="200" swimtime="00:02:02.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196794" lastname="PIGREE" firstname="Analia" gender="F" birthdate="2001-07-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.40" eventid="2" heat="5" lane="3">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.96" eventid="18" heat="6" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="24" lane="3" heat="5" heatid="50002" swimtime="00:00:58.50" reactiontime="+54" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:43.43" />
                    <SPLIT distance="100" swimtime="00:00:58.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="16" lane="5" heat="6" heatid="60018" swimtime="00:00:26.54" reactiontime="+55" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="11" lane="8" heat="1" heatid="10218" swimtime="00:00:26.26" reactiontime="+54" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100908" lastname="BONNET" firstname="Charlotte" gender="F" birthdate="1995-02-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.03" eventid="15" heat="5" lane="2">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.34" eventid="28" heat="3" lane="2">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.69" eventid="6" heat="3" lane="6">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:30.06" eventid="40" heat="7" lane="7">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="15" lane="2" heat="5" heatid="50015" swimtime="00:01:05.28" reactiontime="+71" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="75" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="16" lane="8" heat="2" heatid="20215" swimtime="00:01:05.51" reactiontime="+71" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="75" swimtime="00:00:48.09" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="15" lane="2" heat="3" heatid="30028" swimtime="00:02:21.94" reactiontime="+67" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="75" swimtime="00:00:49.64" />
                    <SPLIT distance="100" swimtime="00:01:07.62" />
                    <SPLIT distance="125" swimtime="00:01:25.89" />
                    <SPLIT distance="150" swimtime="00:01:44.57" />
                    <SPLIT distance="175" swimtime="00:02:03.29" />
                    <SPLIT distance="200" swimtime="00:02:21.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106" place="7" lane="2" heat="1" heatid="10106" swimtime="00:02:07.37" reactiontime="+71" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.25" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:00.10" />
                    <SPLIT distance="125" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:01:37.39" />
                    <SPLIT distance="175" swimtime="00:01:53.34" />
                    <SPLIT distance="200" swimtime="00:02:07.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="5" lane="6" heat="3" heatid="30006" swimtime="00:02:06.70" reactiontime="+71" points="889">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="75" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:00:59.58" />
                    <SPLIT distance="125" swimtime="00:01:18.08" />
                    <SPLIT distance="150" swimtime="00:01:36.64" />
                    <SPLIT distance="175" swimtime="00:01:52.53" />
                    <SPLIT distance="200" swimtime="00:02:06.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="17" lane="7" heat="7" heatid="70040" swimtime="00:00:30.35" reactiontime="+68" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.90" />
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121265" lastname="GASTALDELLO" firstname="Beryl " gender="F" birthdate="1995-02-16">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:51.67" eventid="13" heat="8" lane="5">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:25.16" eventid="4" heat="4" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:00:57.76" eventid="22" heat="4" lane="4">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="7" lane="2" heat="1" heatid="10113" swimtime="00:00:52.13" reactiontime="+64" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:24.83" />
                    <SPLIT distance="75" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:00:52.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="4" lane="5" heat="8" heatid="80013" swimtime="00:00:52.34" reactiontime="+64" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="75" swimtime="00:00:38.60" />
                    <SPLIT distance="100" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="5" lane="5" heat="1" heatid="10213" swimtime="00:00:52.09" reactiontime="+64" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:24.79" />
                    <SPLIT distance="75" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:00:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="104" place="4" lane="1" heat="1" heatid="10104" swimtime="00:00:24.85" reactiontime="+66" points="944">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:24.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="7" lane="3" heat="4" heatid="40004" swimtime="00:00:25.30" reactiontime="+64" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.52" />
                    <SPLIT distance="50" swimtime="00:00:25.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="7" lane="6" heat="2" heatid="20204" swimtime="00:00:25.06" reactiontime="+63" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:25.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="2" lane="6" heat="1" heatid="10122" swimtime="00:00:57.63" reactiontime="+63" points="942">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="75" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:00:57.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="5" lane="4" heat="4" heatid="40022" swimtime="00:00:59.19" reactiontime="+64" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="75" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:00:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="4" lane="3" heat="1" heatid="10222" swimtime="00:00:58.61" reactiontime="+64" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                    <SPLIT distance="75" swimtime="00:00:44.27" />
                    <SPLIT distance="100" swimtime="00:00:58.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129474" lastname="TEREBO" firstname="Emma" gender="F" birthdate="1998-07-10">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.28" eventid="45" heat="3" lane="7">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="17" lane="7" heat="3" heatid="30045" swimtime="00:02:05.94" reactiontime="+57" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="75" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:01.24" />
                    <SPLIT distance="125" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:01:33.86" />
                    <SPLIT distance="175" swimtime="00:01:50.20" />
                    <SPLIT distance="200" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129283" lastname="DUHAMEL" firstname="Cyrielle" gender="F" birthdate="2000-01-06">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.84" eventid="6" heat="3" lane="1">
                  <MEETINFO date="2021-07-27" />
                </ENTRY>
                <ENTRY entrytime="00:04:33.82" eventid="36" heat="4" lane="1">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="23" lane="1" heat="3" heatid="30006" swimtime="00:02:11.20" reactiontime="+67" points="801">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="75" swimtime="00:00:46.29" />
                    <SPLIT distance="100" swimtime="00:01:03.04" />
                    <SPLIT distance="125" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:01:40.51" />
                    <SPLIT distance="175" swimtime="00:01:56.63" />
                    <SPLIT distance="200" swimtime="00:02:11.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="6" lane="8" heat="1" heatid="10136" swimtime="00:04:32.40" reactiontime="+66" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                    <SPLIT distance="75" swimtime="00:00:45.16" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                    <SPLIT distance="125" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:01:37.17" />
                    <SPLIT distance="175" swimtime="00:01:54.46" />
                    <SPLIT distance="200" swimtime="00:02:11.53" />
                    <SPLIT distance="225" swimtime="00:02:30.93" />
                    <SPLIT distance="250" swimtime="00:02:50.20" />
                    <SPLIT distance="275" swimtime="00:03:09.76" />
                    <SPLIT distance="300" swimtime="00:03:29.42" />
                    <SPLIT distance="325" swimtime="00:03:45.58" />
                    <SPLIT distance="350" swimtime="00:04:01.29" />
                    <SPLIT distance="375" swimtime="00:04:17.07" />
                    <SPLIT distance="400" swimtime="00:04:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="8" lane="1" heat="4" heatid="40036" swimtime="00:04:34.03" reactiontime="+66" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.02" />
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="75" swimtime="00:00:45.36" />
                    <SPLIT distance="100" swimtime="00:01:01.97" />
                    <SPLIT distance="125" swimtime="00:01:20.23" />
                    <SPLIT distance="150" swimtime="00:01:37.72" />
                    <SPLIT distance="175" swimtime="00:01:55.26" />
                    <SPLIT distance="200" swimtime="00:02:12.76" />
                    <SPLIT distance="225" swimtime="00:02:31.92" />
                    <SPLIT distance="250" swimtime="00:02:51.44" />
                    <SPLIT distance="275" swimtime="00:03:10.88" />
                    <SPLIT distance="300" swimtime="00:03:30.65" />
                    <SPLIT distance="325" swimtime="00:03:46.84" />
                    <SPLIT distance="350" swimtime="00:04:02.63" />
                    <SPLIT distance="375" swimtime="00:04:18.52" />
                    <SPLIT distance="400" swimtime="00:04:34.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210294" lastname="REYNA" firstname="Alexa" gender="F" birthdate="2005-10-25">
              <ENTRIES>
                <ENTRY entrytime="00:04:06.93" eventid="1" heat="2" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:08:29.84" eventid="12" heat="2" lane="2">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:16:02.61" eventid="33" heat="0" lane="2147483647">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="14" lane="4" heat="2" heatid="20001" swimtime="00:04:08.44" reactiontime="+70" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                    <SPLIT distance="75" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:00:59.35" />
                    <SPLIT distance="125" swimtime="00:01:15.05" />
                    <SPLIT distance="150" swimtime="00:01:30.78" />
                    <SPLIT distance="175" swimtime="00:01:46.58" />
                    <SPLIT distance="200" swimtime="00:02:02.34" />
                    <SPLIT distance="225" swimtime="00:02:18.23" />
                    <SPLIT distance="250" swimtime="00:02:33.95" />
                    <SPLIT distance="275" swimtime="00:02:49.94" />
                    <SPLIT distance="300" swimtime="00:03:05.88" />
                    <SPLIT distance="325" swimtime="00:03:21.73" />
                    <SPLIT distance="350" swimtime="00:03:37.47" />
                    <SPLIT distance="375" swimtime="00:03:53.28" />
                    <SPLIT distance="400" swimtime="00:04:08.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="12" lane="2" heat="2" heatid="20012" swimtime="00:08:35.32" reactiontime="+70" points="804">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="75" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:00.43" />
                    <SPLIT distance="125" swimtime="00:01:16.33" />
                    <SPLIT distance="150" swimtime="00:01:32.26" />
                    <SPLIT distance="175" swimtime="00:01:48.33" />
                    <SPLIT distance="200" swimtime="00:02:04.40" />
                    <SPLIT distance="225" swimtime="00:02:20.32" />
                    <SPLIT distance="250" swimtime="00:02:36.32" />
                    <SPLIT distance="275" swimtime="00:02:52.34" />
                    <SPLIT distance="300" swimtime="00:03:08.42" />
                    <SPLIT distance="325" swimtime="00:03:24.49" />
                    <SPLIT distance="350" swimtime="00:03:40.69" />
                    <SPLIT distance="375" swimtime="00:03:56.79" />
                    <SPLIT distance="400" swimtime="00:04:12.91" />
                    <SPLIT distance="425" swimtime="00:04:28.99" />
                    <SPLIT distance="450" swimtime="00:04:45.28" />
                    <SPLIT distance="475" swimtime="00:05:01.44" />
                    <SPLIT distance="500" swimtime="00:05:17.80" />
                    <SPLIT distance="525" swimtime="00:05:34.08" />
                    <SPLIT distance="550" swimtime="00:05:50.46" />
                    <SPLIT distance="575" swimtime="00:06:06.87" />
                    <SPLIT distance="600" swimtime="00:06:23.25" />
                    <SPLIT distance="625" swimtime="00:06:39.72" />
                    <SPLIT distance="650" swimtime="00:06:56.46" />
                    <SPLIT distance="675" swimtime="00:07:13.02" />
                    <SPLIT distance="700" swimtime="00:07:29.62" />
                    <SPLIT distance="725" swimtime="00:07:46.25" />
                    <SPLIT distance="750" swimtime="00:08:02.83" />
                    <SPLIT distance="775" swimtime="00:08:19.35" />
                    <SPLIT distance="800" swimtime="00:08:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="11" lane="7" heat="5" heatid="30133" swimtime="00:16:23.32" reactiontime="+71" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.89" />
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="75" swimtime="00:00:45.11" />
                    <SPLIT distance="100" swimtime="00:01:00.98" />
                    <SPLIT distance="125" swimtime="00:01:16.95" />
                    <SPLIT distance="150" swimtime="00:01:32.88" />
                    <SPLIT distance="175" swimtime="00:01:48.76" />
                    <SPLIT distance="200" swimtime="00:02:04.70" />
                    <SPLIT distance="225" swimtime="00:02:20.69" />
                    <SPLIT distance="250" swimtime="00:02:36.70" />
                    <SPLIT distance="275" swimtime="00:02:52.69" />
                    <SPLIT distance="300" swimtime="00:03:08.74" />
                    <SPLIT distance="325" swimtime="00:03:24.87" />
                    <SPLIT distance="350" swimtime="00:03:41.00" />
                    <SPLIT distance="375" swimtime="00:03:57.10" />
                    <SPLIT distance="400" swimtime="00:04:13.34" />
                    <SPLIT distance="425" swimtime="00:04:29.53" />
                    <SPLIT distance="450" swimtime="00:04:45.89" />
                    <SPLIT distance="475" swimtime="00:05:02.25" />
                    <SPLIT distance="500" swimtime="00:05:18.71" />
                    <SPLIT distance="525" swimtime="00:05:35.01" />
                    <SPLIT distance="550" swimtime="00:05:51.52" />
                    <SPLIT distance="575" swimtime="00:06:07.91" />
                    <SPLIT distance="600" swimtime="00:06:24.39" />
                    <SPLIT distance="625" swimtime="00:06:40.90" />
                    <SPLIT distance="650" swimtime="00:06:57.56" />
                    <SPLIT distance="675" swimtime="00:07:14.12" />
                    <SPLIT distance="700" swimtime="00:07:30.75" />
                    <SPLIT distance="725" swimtime="00:07:47.23" />
                    <SPLIT distance="750" swimtime="00:08:03.79" />
                    <SPLIT distance="775" swimtime="00:08:20.24" />
                    <SPLIT distance="800" swimtime="00:08:37.03" />
                    <SPLIT distance="825" swimtime="00:08:53.49" />
                    <SPLIT distance="850" swimtime="00:09:10.22" />
                    <SPLIT distance="875" swimtime="00:09:26.83" />
                    <SPLIT distance="900" swimtime="00:09:43.42" />
                    <SPLIT distance="925" swimtime="00:09:59.97" />
                    <SPLIT distance="950" swimtime="00:10:16.67" />
                    <SPLIT distance="975" swimtime="00:10:33.15" />
                    <SPLIT distance="1000" swimtime="00:10:49.90" />
                    <SPLIT distance="1025" swimtime="00:11:06.52" />
                    <SPLIT distance="1050" swimtime="00:11:23.32" />
                    <SPLIT distance="1075" swimtime="00:11:39.97" />
                    <SPLIT distance="1100" swimtime="00:11:56.64" />
                    <SPLIT distance="1125" swimtime="00:12:13.36" />
                    <SPLIT distance="1150" swimtime="00:12:30.23" />
                    <SPLIT distance="1175" swimtime="00:12:47.00" />
                    <SPLIT distance="1200" swimtime="00:13:03.82" />
                    <SPLIT distance="1225" swimtime="00:13:20.52" />
                    <SPLIT distance="1250" swimtime="00:13:37.30" />
                    <SPLIT distance="1275" swimtime="00:13:53.91" />
                    <SPLIT distance="1300" swimtime="00:14:10.71" />
                    <SPLIT distance="1325" swimtime="00:14:27.47" />
                    <SPLIT distance="1350" swimtime="00:14:44.20" />
                    <SPLIT distance="1375" swimtime="00:15:00.76" />
                    <SPLIT distance="1400" swimtime="00:15:17.48" />
                    <SPLIT distance="1425" swimtime="00:15:33.98" />
                    <SPLIT distance="1450" swimtime="00:15:50.49" />
                    <SPLIT distance="1475" swimtime="00:16:06.98" />
                    <SPLIT distance="1500" swimtime="00:16:23.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197599" lastname="MOLUH" firstname="Mary-Ambre" gender="F" birthdate="2005-09-09">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:26.33" eventid="18" heat="5" lane="6">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="14" lane="6" heat="5" heatid="50018" swimtime="00:00:26.45" reactiontime="+62" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="15" lane="1" heat="1" heatid="10218" swimtime="00:00:26.54" reactiontime="+61" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100470" lastname="HENIQUE" firstname="Melanie" gender="F" birthdate="1992-12-22">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:24.91" eventid="4" heat="5" lane="5">
                  <MEETINFO date="2021-11-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.95" eventid="30" heat="7" lane="6">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="104" place="5" lane="2" heat="1" heatid="10104" swimtime="00:00:24.92" reactiontime="+59" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.18" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="2" lane="5" heat="5" heatid="50004" swimtime="00:00:24.88" reactiontime="+58" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.07" />
                    <SPLIT distance="50" swimtime="00:00:24.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="4" lane="4" heat="1" heatid="10204" swimtime="00:00:24.92" reactiontime="+57" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="8" lane="8" heat="1" heatid="10130" swimtime="00:00:23.90" reactiontime="+59" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:23.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="4" lane="6" heat="7" heatid="70030" swimtime="00:00:23.86" reactiontime="+59" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:23.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="7" lane="3" heat="2" heatid="20230" swimtime="00:00:24.00" reactiontime="+57" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:24.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121517" lastname="BOUCHAUT" firstname="Joris " gender="M" birthdate="1995-06-27">
              <ENTRIES>
                <ENTRY entrytime="00:07:36.22" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="142" place="6" lane="6" heat="5" heatid="30142" swimtime="00:07:35.12" reactiontime="+72" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                    <SPLIT distance="75" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:00:55.12" />
                    <SPLIT distance="125" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:23.66" />
                    <SPLIT distance="175" swimtime="00:01:37.74" />
                    <SPLIT distance="200" swimtime="00:01:51.97" />
                    <SPLIT distance="225" swimtime="00:02:06.14" />
                    <SPLIT distance="250" swimtime="00:02:20.40" />
                    <SPLIT distance="275" swimtime="00:02:34.74" />
                    <SPLIT distance="300" swimtime="00:02:49.21" />
                    <SPLIT distance="325" swimtime="00:03:03.55" />
                    <SPLIT distance="350" swimtime="00:03:17.86" />
                    <SPLIT distance="375" swimtime="00:03:32.41" />
                    <SPLIT distance="400" swimtime="00:03:46.74" />
                    <SPLIT distance="425" swimtime="00:04:00.92" />
                    <SPLIT distance="450" swimtime="00:04:15.28" />
                    <SPLIT distance="475" swimtime="00:04:29.23" />
                    <SPLIT distance="500" swimtime="00:04:43.47" />
                    <SPLIT distance="525" swimtime="00:04:57.53" />
                    <SPLIT distance="550" swimtime="00:05:11.71" />
                    <SPLIT distance="575" swimtime="00:05:25.94" />
                    <SPLIT distance="600" swimtime="00:05:40.24" />
                    <SPLIT distance="625" swimtime="00:05:54.59" />
                    <SPLIT distance="650" swimtime="00:06:09.05" />
                    <SPLIT distance="675" swimtime="00:06:23.57" />
                    <SPLIT distance="700" swimtime="00:06:38.19" />
                    <SPLIT distance="725" swimtime="00:06:52.64" />
                    <SPLIT distance="750" swimtime="00:07:07.41" />
                    <SPLIT distance="775" swimtime="00:07:21.70" />
                    <SPLIT distance="800" swimtime="00:07:35.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="France">
              <RESULTS>
                <RESULT eventid="127" place="1" lane="4" heat="1" swimtime="00:01:27.33" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.13" />
                    <SPLIT distance="50" swimtime="00:00:20.92" />
                    <SPLIT distance="75" swimtime="00:00:30.32" />
                    <SPLIT distance="100" swimtime="00:00:41.18" />
                    <SPLIT distance="125" swimtime="00:00:51.85" />
                    <SPLIT distance="150" swimtime="00:01:04.18" />
                    <SPLIT distance="175" swimtime="00:01:14.95" />
                    <SPLIT distance="200" swimtime="00:01:27.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="149769" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="101299" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="121265" reactiontime="+9" />
                    <RELAYPOSITION number="4" athleteid="100470" reactiontime="+1" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="1" lane="5" heat="3" swimtime="00:01:29.69" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.16" />
                    <SPLIT distance="50" swimtime="00:00:21.10" />
                    <SPLIT distance="75" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:00:41.86" />
                    <SPLIT distance="125" swimtime="00:00:53.03" />
                    <SPLIT distance="150" swimtime="00:01:05.72" />
                    <SPLIT distance="175" swimtime="00:01:17.15" />
                    <SPLIT distance="200" swimtime="00:01:29.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101299" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="149769" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="100470" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="197599" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="France">
              <RESULTS>
                <RESULT eventid="147" place="6" lane="1" heat="1" swimtime="00:03:50.28" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="75" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:00:57.22" />
                    <SPLIT distance="125" swimtime="00:01:10.66" />
                    <SPLIT distance="150" swimtime="00:01:27.20" />
                    <SPLIT distance="175" swimtime="00:01:44.07" />
                    <SPLIT distance="200" swimtime="00:02:01.34" />
                    <SPLIT distance="225" swimtime="00:02:12.76" />
                    <SPLIT distance="250" swimtime="00:02:26.83" />
                    <SPLIT distance="275" swimtime="00:02:41.92" />
                    <SPLIT distance="300" swimtime="00:02:57.54" />
                    <SPLIT distance="325" swimtime="00:03:09.24" />
                    <SPLIT distance="350" swimtime="00:03:22.53" />
                    <SPLIT distance="375" swimtime="00:03:36.35" />
                    <SPLIT distance="400" swimtime="00:03:50.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="110511" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="100908" reactiontime="+12" />
                    <RELAYPOSITION number="3" athleteid="121265" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="197599" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="7" lane="6" heat="1" swimtime="00:03:53.55" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="75" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:00:57.36" />
                    <SPLIT distance="125" swimtime="00:01:11.42" />
                    <SPLIT distance="150" swimtime="00:01:28.39" />
                    <SPLIT distance="175" swimtime="00:01:45.69" />
                    <SPLIT distance="200" swimtime="00:02:02.94" />
                    <SPLIT distance="225" swimtime="00:02:14.57" />
                    <SPLIT distance="250" swimtime="00:02:28.93" />
                    <SPLIT distance="275" swimtime="00:02:43.93" />
                    <SPLIT distance="300" swimtime="00:02:59.84" />
                    <SPLIT distance="325" swimtime="00:03:11.15" />
                    <SPLIT distance="350" swimtime="00:03:24.44" />
                    <SPLIT distance="375" swimtime="00:03:38.76" />
                    <SPLIT distance="400" swimtime="00:03:53.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197599" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="100908" reactiontime="+30" />
                    <RELAYPOSITION number="3" athleteid="121265" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="100470" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="France">
              <RESULTS>
                <RESULT eventid="134" place="6" lane="3" heat="1" swimtime="00:01:43.96" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.96" />
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                    <SPLIT distance="75" swimtime="00:00:39.80" />
                    <SPLIT distance="100" swimtime="00:00:55.94" />
                    <SPLIT distance="125" swimtime="00:01:07.05" />
                    <SPLIT distance="150" swimtime="00:01:20.72" />
                    <SPLIT distance="175" swimtime="00:01:31.73" />
                    <SPLIT distance="200" swimtime="00:01:43.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196794" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="100908" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="100470" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="121265" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="3" lane="6" heat="2" swimtime="00:01:44.86" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.06" />
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="75" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:00:56.12" />
                    <SPLIT distance="125" swimtime="00:01:07.50" />
                    <SPLIT distance="150" swimtime="00:01:21.48" />
                    <SPLIT distance="175" swimtime="00:01:32.48" />
                    <SPLIT distance="200" swimtime="00:01:44.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196794" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="100908" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="100470" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="121265" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="France">
              <RESULTS>
                <RESULT eventid="135" place="5" lane="5" heat="1" swimtime="00:01:31.41" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.30" />
                    <SPLIT distance="50" swimtime="00:00:22.96" />
                    <SPLIT distance="75" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:00:48.97" />
                    <SPLIT distance="125" swimtime="00:00:58.74" />
                    <SPLIT distance="150" swimtime="00:01:10.87" />
                    <SPLIT distance="175" swimtime="00:01:20.44" />
                    <SPLIT distance="200" swimtime="00:01:31.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="181969" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="201991" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="149769" reactiontime="+7" />
                    <RELAYPOSITION number="4" athleteid="101299" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="2" lane="7" heat="3" swimtime="00:01:32.53" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:23.44" />
                    <SPLIT distance="75" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:00:49.62" />
                    <SPLIT distance="125" swimtime="00:00:59.70" />
                    <SPLIT distance="150" swimtime="00:01:11.80" />
                    <SPLIT distance="175" swimtime="00:01:21.52" />
                    <SPLIT distance="200" swimtime="00:01:32.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="191730" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="197601" reactiontime="+45" />
                    <RELAYPOSITION number="3" athleteid="149769" reactiontime="+40" />
                    <RELAYPOSITION number="4" athleteid="101299" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="" shortname="FRO" code="FRO" nation="" type="">
          <ATHLETES>
            <ATHLETE athleteid="125170" lastname="EIDESGAARD" firstname="Var" gender="F" birthdate="2001-03-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.60" eventid="13" heat="4" lane="4">
                  <MEETINFO date="2022-11-11" />
                </ENTRY>
                <ENTRY entrytime="00:04:14.09" eventid="1" heat="2" lane="8">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="40" lane="4" heat="4" heatid="40013" swimtime="00:00:56.21" reactiontime="+66" points="714">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="75" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:00:56.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="22" lane="8" heat="2" heatid="20001" swimtime="00:04:16.97" reactiontime="+70" points="754">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.85" />
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="75" swimtime="00:00:45.26" />
                    <SPLIT distance="100" swimtime="00:01:01.18" />
                    <SPLIT distance="125" swimtime="00:01:17.43" />
                    <SPLIT distance="150" swimtime="00:01:33.53" />
                    <SPLIT distance="175" swimtime="00:01:49.90" />
                    <SPLIT distance="200" swimtime="00:02:06.29" />
                    <SPLIT distance="225" swimtime="00:02:22.70" />
                    <SPLIT distance="250" swimtime="00:02:39.12" />
                    <SPLIT distance="275" swimtime="00:02:55.82" />
                    <SPLIT distance="300" swimtime="00:03:12.22" />
                    <SPLIT distance="325" swimtime="00:03:28.74" />
                    <SPLIT distance="350" swimtime="00:03:45.15" />
                    <SPLIT distance="375" swimtime="00:04:01.63" />
                    <SPLIT distance="400" swimtime="00:04:16.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Micronesia" shortname="FSM" code="FSM" nation="FSM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154951" lastname="LIMTIACO" firstname="Tasi" gender="M" birthdate="1994-01-04">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.16" eventid="16" heat="2" lane="2">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.23" eventid="41" heat="3" lane="6">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="52" lane="2" heat="2" heatid="20016" swimtime="00:01:01.98" reactiontime="+66" points="709">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                    <SPLIT distance="75" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="45" lane="6" heat="3" heatid="30041" swimtime="00:00:28.26" reactiontime="+68" points="688">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201593" lastname="KIHLENG" firstname="Kyler Anthony" gender="M" birthdate="2004-12-23">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.95" eventid="14" heat="2" lane="8">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.95" eventid="31" heat="3" lane="7">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="82" lane="8" heat="2" heatid="20014" swimtime="00:00:58.58" reactiontime="+69" points="448">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                    <SPLIT distance="75" swimtime="00:00:43.66" />
                    <SPLIT distance="100" swimtime="00:00:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="69" lane="7" heat="3" heatid="30031" swimtime="00:00:26.47" reactiontime="+66" points="441">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130104" lastname="ADAMS" firstname="Taeyanna" gender="F" birthdate="2002-03-14">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:36.11" eventid="40" heat="3" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="37" lane="8" heat="3" heatid="30040" swimtime="00:00:36.64" reactiontime="+69" points="473">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="45" lane="4" heat="1" heatid="10030" swimtime="00:00:28.84" reactiontime="+66" points="502">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130130" lastname="KIHLENG" firstname="Kestra" gender="F" birthdate="2003-08-12">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:31.76" eventid="4" heat="2" lane="2">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="6" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="37" lane="2" heat="2" heatid="20004" swimtime="00:00:31.25" reactiontime="+70" points="474">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="29" lane="6" heat="1" heatid="10022" swimtime="00:01:14.77" reactiontime="+66" points="431">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                    <SPLIT distance="75" swimtime="00:00:55.91" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Federated States of Micronesia">
              <RESULTS>
                <RESULT eventid="27" place="25" lane="1" heat="4" swimtime="00:01:48.53" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                    <SPLIT distance="75" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:00:53.32" />
                    <SPLIT distance="125" swimtime="00:01:07.17" />
                    <SPLIT distance="150" swimtime="00:01:22.51" />
                    <SPLIT distance="175" swimtime="00:01:35.13" />
                    <SPLIT distance="200" swimtime="00:01:48.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154951" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="130104" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="130130" reactiontime="+14" />
                    <RELAYPOSITION number="4" athleteid="201593" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Federated States of Micronesia">
              <RESULTS>
                <RESULT eventid="11" place="29" lane="3" heat="1" swimtime="00:02:02.75" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                    <SPLIT distance="75" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:04.69" />
                    <SPLIT distance="125" swimtime="00:01:18.79" />
                    <SPLIT distance="150" swimtime="00:01:36.29" />
                    <SPLIT distance="175" swimtime="00:01:49.37" />
                    <SPLIT distance="200" swimtime="00:02:02.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154951" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="130104" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="130130" reactiontime="+17" />
                    <RELAYPOSITION number="4" athleteid="201593" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Gambia" shortname="GAM" code="GAM" nation="GAM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="110890" lastname="JONGA" firstname="Pap D" gender="M" birthdate="1997-07-01">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="31" heat="1" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="64" lane="3" heat="1" heatid="10005" swimtime="00:00:29.20" reactiontime="+77" points="413">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="72" lane="6" heat="1" heatid="10031" swimtime="00:00:26.73" reactiontime="+69" points="429">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Great Britain" shortname="GBR" code="GBR" nation="GBR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="125048" lastname="GREENBANK" firstname="Luke" gender="M" birthdate="1997-09-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.48" eventid="3" heat="4" lane="3">
                  <MEETINFO date="2021-09-02" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.15" eventid="46" heat="3" lane="3">
                  <MEETINFO date="2021-09-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="13" lane="3" heat="4" heatid="40003" swimtime="00:00:50.72" reactiontime="+57" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.81" />
                    <SPLIT distance="50" swimtime="00:00:24.42" />
                    <SPLIT distance="75" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:00:50.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="14" lane="1" heat="2" heatid="20203" swimtime="00:00:50.81" reactiontime="+56" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:24.76" />
                    <SPLIT distance="75" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="146" place="5" lane="7" heat="1" heatid="10146" swimtime="00:01:49.79" reactiontime="+60" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:26.19" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:54.27" />
                    <SPLIT distance="125" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:22.12" />
                    <SPLIT distance="175" swimtime="00:01:36.09" />
                    <SPLIT distance="200" swimtime="00:01:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="6" lane="3" heat="3" heatid="30046" swimtime="00:01:50.34" reactiontime="+60" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:00:53.48" />
                    <SPLIT distance="125" swimtime="00:01:07.62" />
                    <SPLIT distance="150" swimtime="00:01:21.69" />
                    <SPLIT distance="175" swimtime="00:01:36.08" />
                    <SPLIT distance="200" swimtime="00:01:50.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108588" lastname="PEATY" firstname="Adam" gender="M" birthdate="1994-12-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.37" eventid="16" heat="7" lane="2">
                  <MEETINFO date="2021-07-26" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.48" eventid="29" heat="1" lane="4">
                  <MEETINFO date="2022-03-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.65" eventid="41" heat="8" lane="1">
                  <MEETINFO date="2021-07-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="3" lane="6" heat="1" heatid="10116" swimtime="00:00:56.25" reactiontime="+61" points="949">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                    <SPLIT distance="75" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:00:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="4" lane="2" heat="7" heatid="70016" swimtime="00:00:56.81" reactiontime="+59" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:26.46" />
                    <SPLIT distance="75" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:00:56.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="4" lane="5" heat="1" heatid="10216" swimtime="00:00:56.42" reactiontime="+58" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:26.41" />
                    <SPLIT distance="75" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:00:56.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="18" lane="4" heat="1" heatid="10029" swimtime="00:02:07.31" reactiontime="+62" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                    <SPLIT distance="75" swimtime="00:00:43.42" />
                    <SPLIT distance="100" swimtime="00:00:59.61" />
                    <SPLIT distance="125" swimtime="00:01:16.00" />
                    <SPLIT distance="150" swimtime="00:01:32.88" />
                    <SPLIT distance="175" swimtime="00:01:49.78" />
                    <SPLIT distance="200" swimtime="00:02:07.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="6" lane="1" heat="1" heatid="10141" swimtime="00:00:25.99" reactiontime="+57" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="2" lane="1" heat="8" heatid="80041" swimtime="00:00:26.01" reactiontime="+60" points="882">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.79" />
                    <SPLIT distance="50" swimtime="00:00:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="7" lane="4" heat="1" heatid="10241" swimtime="00:00:25.85" reactiontime="+61" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150500" lastname="BURRAS" firstname="Lewis Edward" gender="M" birthdate="2000-02-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.63" eventid="14" heat="8" lane="6">
                  <MEETINFO date="2022-06-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.55" eventid="5" heat="5" lane="3">
                  <MEETINFO date="2022-05-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.68" eventid="31" heat="8" lane="2">
                  <MEETINFO date="2022-08-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="13" lane="6" heat="8" heatid="80014" swimtime="00:00:46.92" reactiontime="+64" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.40" />
                    <SPLIT distance="50" swimtime="00:00:22.05" />
                    <SPLIT distance="75" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:00:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="12" lane="1" heat="2" heatid="20214" swimtime="00:00:46.61" reactiontime="+61" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.37" />
                    <SPLIT distance="50" swimtime="00:00:22.11" />
                    <SPLIT distance="75" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:00:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="35" lane="3" heat="5" heatid="50005" swimtime="00:00:23.18" reactiontime="+64" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="131" place="8" lane="2" heat="1" heatid="10131" swimtime="00:00:20.95" reactiontime="+60" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.13" />
                    <SPLIT distance="50" swimtime="00:00:20.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="6" lane="2" heat="8" heatid="80031" swimtime="00:00:21.00" reactiontime="+61" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.16" />
                    <SPLIT distance="50" swimtime="00:00:21.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="5" lane="3" heat="1" heatid="10231" swimtime="00:00:20.94" reactiontime="+65" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.22" />
                    <SPLIT distance="50" swimtime="00:00:20.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165917" lastname="DEAN" firstname="Tom" gender="M" birthdate="2000-05-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.83" eventid="14" heat="8" lane="2">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.25" eventid="44" heat="5" lane="7">
                  <MEETINFO date="2021-12-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:56.77" eventid="7" heat="4" lane="1">
                  <MEETINFO date="2022-06-22" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.20" eventid="24" heat="5" lane="1">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="8" lane="8" heat="1" heatid="10114" swimtime="00:00:46.11" reactiontime="+70" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.55" />
                    <SPLIT distance="50" swimtime="00:00:22.16" />
                    <SPLIT distance="75" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="9" lane="2" heat="8" heatid="80014" swimtime="00:00:46.54" reactiontime="+67" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.57" />
                    <SPLIT distance="50" swimtime="00:00:22.23" />
                    <SPLIT distance="75" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="8" lane="2" heat="2" heatid="20214" swimtime="00:00:46.20" reactiontime="+65" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.53" />
                    <SPLIT distance="50" swimtime="00:00:22.15" />
                    <SPLIT distance="75" swimtime="00:00:34.22" />
                    <SPLIT distance="100" swimtime="00:00:46.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="144" place="3" lane="4" heat="1" heatid="10144" swimtime="00:01:40.86" reactiontime="+65" points="956">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.99" />
                    <SPLIT distance="50" swimtime="00:00:23.35" />
                    <SPLIT distance="75" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:00:48.81" />
                    <SPLIT distance="125" swimtime="00:01:01.82" />
                    <SPLIT distance="150" swimtime="00:01:15.09" />
                    <SPLIT distance="175" swimtime="00:01:28.14" />
                    <SPLIT distance="200" swimtime="00:01:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="1" lane="7" heat="5" heatid="50044" swimtime="00:01:40.98" reactiontime="+66" points="952">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.92" />
                    <SPLIT distance="50" swimtime="00:00:23.20" />
                    <SPLIT distance="75" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:00:48.64" />
                    <SPLIT distance="125" swimtime="00:01:01.53" />
                    <SPLIT distance="150" swimtime="00:01:14.82" />
                    <SPLIT distance="175" swimtime="00:01:28.19" />
                    <SPLIT distance="200" swimtime="00:01:40.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="11" lane="1" heat="4" heatid="40007" swimtime="00:01:53.53" reactiontime="+71" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.88" />
                    <SPLIT distance="50" swimtime="00:00:24.36" />
                    <SPLIT distance="75" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:00:52.93" />
                    <SPLIT distance="125" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:26.17" />
                    <SPLIT distance="175" swimtime="00:01:40.65" />
                    <SPLIT distance="200" swimtime="00:01:53.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="10" lane="1" heat="5" heatid="50024" swimtime="00:03:39.79" reactiontime="+68" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                    <SPLIT distance="75" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:00:51.65" />
                    <SPLIT distance="125" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:19.48" />
                    <SPLIT distance="175" swimtime="00:01:33.31" />
                    <SPLIT distance="200" swimtime="00:01:47.41" />
                    <SPLIT distance="225" swimtime="00:02:01.29" />
                    <SPLIT distance="250" swimtime="00:02:15.37" />
                    <SPLIT distance="275" swimtime="00:02:29.33" />
                    <SPLIT distance="300" swimtime="00:02:43.55" />
                    <SPLIT distance="325" swimtime="00:02:57.70" />
                    <SPLIT distance="350" swimtime="00:03:11.99" />
                    <SPLIT distance="375" swimtime="00:03:26.22" />
                    <SPLIT distance="400" swimtime="00:03:39.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144828" lastname="JERVIS" firstname="Daniel" gender="M" birthdate="1996-06-09">
              <ENTRIES>
                <ENTRY entrytime="00:14:48.86" eventid="10" heat="2" lane="7">
                  <MEETINFO date="2022-06-25" />
                </ENTRY>
                <ENTRY entrytime="00:03:46.44" eventid="24" heat="3" lane="1">
                  <MEETINFO date="2022-04-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="6" lane="7" heat="2" heatid="20010" swimtime="00:14:30.47" reactiontime="+63" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="75" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:00:53.96" />
                    <SPLIT distance="125" swimtime="00:01:08.22" />
                    <SPLIT distance="150" swimtime="00:01:22.61" />
                    <SPLIT distance="175" swimtime="00:01:36.93" />
                    <SPLIT distance="200" swimtime="00:01:51.38" />
                    <SPLIT distance="225" swimtime="00:02:05.74" />
                    <SPLIT distance="250" swimtime="00:02:20.18" />
                    <SPLIT distance="275" swimtime="00:02:34.66" />
                    <SPLIT distance="300" swimtime="00:02:49.18" />
                    <SPLIT distance="325" swimtime="00:03:03.56" />
                    <SPLIT distance="350" swimtime="00:03:18.12" />
                    <SPLIT distance="375" swimtime="00:03:32.59" />
                    <SPLIT distance="400" swimtime="00:03:47.16" />
                    <SPLIT distance="425" swimtime="00:04:01.78" />
                    <SPLIT distance="450" swimtime="00:04:16.52" />
                    <SPLIT distance="475" swimtime="00:04:31.21" />
                    <SPLIT distance="500" swimtime="00:04:45.94" />
                    <SPLIT distance="525" swimtime="00:05:00.56" />
                    <SPLIT distance="550" swimtime="00:05:15.23" />
                    <SPLIT distance="575" swimtime="00:05:29.83" />
                    <SPLIT distance="600" swimtime="00:05:44.71" />
                    <SPLIT distance="625" swimtime="00:05:59.47" />
                    <SPLIT distance="650" swimtime="00:06:14.24" />
                    <SPLIT distance="675" swimtime="00:06:28.86" />
                    <SPLIT distance="700" swimtime="00:06:43.66" />
                    <SPLIT distance="725" swimtime="00:06:58.39" />
                    <SPLIT distance="750" swimtime="00:07:13.25" />
                    <SPLIT distance="775" swimtime="00:07:28.11" />
                    <SPLIT distance="800" swimtime="00:07:42.91" />
                    <SPLIT distance="825" swimtime="00:07:57.65" />
                    <SPLIT distance="850" swimtime="00:08:12.45" />
                    <SPLIT distance="875" swimtime="00:08:27.22" />
                    <SPLIT distance="900" swimtime="00:08:41.90" />
                    <SPLIT distance="925" swimtime="00:08:56.47" />
                    <SPLIT distance="950" swimtime="00:09:11.13" />
                    <SPLIT distance="975" swimtime="00:09:25.59" />
                    <SPLIT distance="1000" swimtime="00:09:40.13" />
                    <SPLIT distance="1025" swimtime="00:09:54.68" />
                    <SPLIT distance="1050" swimtime="00:10:09.17" />
                    <SPLIT distance="1075" swimtime="00:10:23.62" />
                    <SPLIT distance="1100" swimtime="00:10:38.57" />
                    <SPLIT distance="1125" swimtime="00:10:53.10" />
                    <SPLIT distance="1150" swimtime="00:11:07.62" />
                    <SPLIT distance="1175" swimtime="00:11:22.16" />
                    <SPLIT distance="1200" swimtime="00:11:36.84" />
                    <SPLIT distance="1225" swimtime="00:11:51.37" />
                    <SPLIT distance="1250" swimtime="00:12:06.07" />
                    <SPLIT distance="1275" swimtime="00:12:20.79" />
                    <SPLIT distance="1300" swimtime="00:12:35.45" />
                    <SPLIT distance="1325" swimtime="00:12:50.11" />
                    <SPLIT distance="1350" swimtime="00:13:04.77" />
                    <SPLIT distance="1375" swimtime="00:13:19.33" />
                    <SPLIT distance="1400" swimtime="00:13:34.09" />
                    <SPLIT distance="1425" swimtime="00:13:48.60" />
                    <SPLIT distance="1450" swimtime="00:14:02.83" />
                    <SPLIT distance="1475" swimtime="00:14:17.01" />
                    <SPLIT distance="1500" swimtime="00:14:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="15" lane="1" heat="3" heatid="30024" swimtime="00:03:42.85" reactiontime="+62" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:25.63" />
                    <SPLIT distance="75" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:00:53.53" />
                    <SPLIT distance="125" swimtime="00:01:07.64" />
                    <SPLIT distance="150" swimtime="00:01:21.91" />
                    <SPLIT distance="175" swimtime="00:01:36.16" />
                    <SPLIT distance="200" swimtime="00:01:50.43" />
                    <SPLIT distance="225" swimtime="00:02:04.66" />
                    <SPLIT distance="250" swimtime="00:02:19.12" />
                    <SPLIT distance="275" swimtime="00:02:33.38" />
                    <SPLIT distance="300" swimtime="00:02:47.55" />
                    <SPLIT distance="325" swimtime="00:03:01.65" />
                    <SPLIT distance="350" swimtime="00:03:15.73" />
                    <SPLIT distance="375" swimtime="00:03:29.64" />
                    <SPLIT distance="400" swimtime="00:03:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101625" lastname="PROUD" firstname="Benjamin" gender="M" birthdate="1994-09-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:20.40" eventid="31" heat="11" lane="4">
                  <MEETINFO date="2021-12-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="131" place="2" lane="5" heat="1" heatid="10131" swimtime="00:00:20.49" reactiontime="+58" points="952">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.81" />
                    <SPLIT distance="50" swimtime="00:00:20.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="3" lane="4" heat="11" heatid="110031" swimtime="00:00:20.88" reactiontime="+58" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.04" />
                    <SPLIT distance="50" swimtime="00:00:20.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="2" lane="5" heat="2" heatid="20231" swimtime="00:00:20.76" reactiontime="+58" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.93" />
                    <SPLIT distance="50" swimtime="00:00:20.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202246" lastname="HARRIS" firstname="Medi Eira" gender="F" birthdate="2002-09-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.46" eventid="2" heat="3" lane="6">
                  <MEETINFO date="2022-08-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="00:00:27.56" eventid="18" heat="6" lane="8">
                  <MEETINFO date="2022-06-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="14" lane="6" heat="3" heatid="30002" swimtime="00:00:57.51" reactiontime="+64" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="75" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="12" lane="1" heat="1" heatid="10202" swimtime="00:00:57.40" reactiontime="+69" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="75" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:00:57.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="17" lane="8" heat="6" heatid="60018" swimtime="00:00:26.68" reactiontime="+64" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161299" lastname="CLARK" firstname="Imogen Louise" gender="F" birthdate="1999-06-01">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.61" eventid="15" heat="4" lane="4">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:29.32" eventid="40" heat="7" lane="5">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="12" lane="4" heat="4" heatid="40015" swimtime="00:01:05.05" reactiontime="+63" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:05.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="14" lane="7" heat="1" heatid="10215" swimtime="00:01:05.40" reactiontime="+64" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="75" swimtime="00:00:47.30" />
                    <SPLIT distance="100" swimtime="00:01:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="6" lane="2" heat="1" heatid="10140" swimtime="00:00:29.47" reactiontime="+65" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="4" lane="5" heat="7" heatid="70040" swimtime="00:00:29.51" reactiontime="+65" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="5" lane="5" heat="1" heatid="10240" swimtime="00:00:29.30" reactiontime="+64" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.36" />
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165928" lastname="HOPKIN" firstname="Anna" gender="F" birthdate="1996-04-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.99" eventid="13" heat="9" lane="6">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:23.89" eventid="30" heat="7" lane="3">
                  <MEETINFO date="2021-11-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="14" lane="6" heat="9" heatid="90013" swimtime="00:00:53.06" reactiontime="+68" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                    <SPLIT distance="75" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:00:53.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="13" lane="1" heat="1" heatid="10213" swimtime="00:00:52.74" reactiontime="+66" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:25.31" />
                    <SPLIT distance="75" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:00:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="3" lane="6" heat="1" heatid="10130" swimtime="00:00:23.68" reactiontime="+67" points="907">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="4" lane="3" heat="7" heatid="70030" swimtime="00:00:23.86" reactiontime="+64" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                    <SPLIT distance="50" swimtime="00:00:23.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="4" lane="5" heat="1" heatid="10230" swimtime="00:00:23.79" reactiontime="+64" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213597" lastname="HINDLEY" firstname="Isabella" gender="F" birthdate="1996-10-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.58" eventid="13" heat="9" lane="2">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:24.20" eventid="30" heat="6" lane="2">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="30" lane="2" heat="9" heatid="90013" swimtime="00:00:54.57" reactiontime="+73" points="780">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="75" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:00:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="19" lane="2" heat="6" heatid="60030" swimtime="00:00:24.86" reactiontime="+70" points="784">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="126805" lastname="WOOD" firstname="Abbie" gender="F" birthdate="1999-03-02">
              <ENTRIES>
                <ENTRY entrytime="00:02:19.11" eventid="28" heat="3" lane="4">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.94" eventid="6" heat="5" lane="5">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:04:27.76" eventid="36" heat="4" lane="5">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="128" place="8" lane="8" heat="1" heatid="10128" swimtime="00:02:21.48" reactiontime="+68" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="75" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                    <SPLIT distance="125" swimtime="00:01:26.00" />
                    <SPLIT distance="150" swimtime="00:01:44.21" />
                    <SPLIT distance="175" swimtime="00:02:02.74" />
                    <SPLIT distance="200" swimtime="00:02:21.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="8" lane="4" heat="3" heatid="30028" swimtime="00:02:20.26" reactiontime="+66" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.64" />
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="75" swimtime="00:00:49.63" />
                    <SPLIT distance="100" swimtime="00:01:07.49" />
                    <SPLIT distance="125" swimtime="00:01:25.60" />
                    <SPLIT distance="150" swimtime="00:01:43.74" />
                    <SPLIT distance="175" swimtime="00:02:02.10" />
                    <SPLIT distance="200" swimtime="00:02:20.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106" place="6" lane="1" heat="1" heatid="10106" swimtime="00:02:07.28" reactiontime="+69" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="75" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:00:59.26" />
                    <SPLIT distance="125" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:01:36.18" />
                    <SPLIT distance="175" swimtime="00:01:52.46" />
                    <SPLIT distance="200" swimtime="00:02:07.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="7" lane="5" heat="5" heatid="50006" swimtime="00:02:07.20" reactiontime="+69" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:27.36" />
                    <SPLIT distance="75" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:00:59.16" />
                    <SPLIT distance="125" swimtime="00:01:17.29" />
                    <SPLIT distance="150" swimtime="00:01:36.19" />
                    <SPLIT distance="175" swimtime="00:01:52.26" />
                    <SPLIT distance="200" swimtime="00:02:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="9" lane="5" heat="4" heatid="40036" swimtime="00:04:34.45" reactiontime="+69" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.23" />
                    <SPLIT distance="50" swimtime="00:00:29.23" />
                    <SPLIT distance="75" swimtime="00:00:45.96" />
                    <SPLIT distance="100" swimtime="00:01:02.85" />
                    <SPLIT distance="125" swimtime="00:01:20.84" />
                    <SPLIT distance="150" swimtime="00:01:38.26" />
                    <SPLIT distance="175" swimtime="00:01:56.01" />
                    <SPLIT distance="200" swimtime="00:02:13.36" />
                    <SPLIT distance="225" swimtime="00:02:32.01" />
                    <SPLIT distance="250" swimtime="00:02:51.08" />
                    <SPLIT distance="275" swimtime="00:03:10.32" />
                    <SPLIT distance="300" swimtime="00:03:29.75" />
                    <SPLIT distance="325" swimtime="00:03:46.57" />
                    <SPLIT distance="350" swimtime="00:04:02.58" />
                    <SPLIT distance="375" swimtime="00:04:18.63" />
                    <SPLIT distance="400" swimtime="00:04:34.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Great Britain">
              <RESULTS>
                <RESULT eventid="48" place="-1" lane="3" heat="2" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Great Britain">
              <RESULTS>
                <RESULT eventid="108" place="7" lane="1" heat="1" swimtime="00:03:33.47" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.79" />
                    <SPLIT distance="50" swimtime="00:00:24.84" />
                    <SPLIT distance="75" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:00:51.81" />
                    <SPLIT distance="125" swimtime="00:01:03.40" />
                    <SPLIT distance="150" swimtime="00:01:17.05" />
                    <SPLIT distance="175" swimtime="00:01:31.18" />
                    <SPLIT distance="200" swimtime="00:01:45.61" />
                    <SPLIT distance="225" swimtime="00:01:58.00" />
                    <SPLIT distance="250" swimtime="00:02:11.70" />
                    <SPLIT distance="275" swimtime="00:02:25.69" />
                    <SPLIT distance="300" swimtime="00:02:39.64" />
                    <SPLIT distance="325" swimtime="00:02:51.64" />
                    <SPLIT distance="350" swimtime="00:03:05.29" />
                    <SPLIT distance="375" swimtime="00:03:19.32" />
                    <SPLIT distance="400" swimtime="00:03:33.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="165928" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="213597" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="202246" reactiontime="+44" />
                    <RELAYPOSITION number="4" athleteid="126805" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="7" lane="6" heat="2" swimtime="00:03:33.46" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:24.76" />
                    <SPLIT distance="75" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:00:52.12" />
                    <SPLIT distance="125" swimtime="00:01:03.83" />
                    <SPLIT distance="150" swimtime="00:01:17.60" />
                    <SPLIT distance="175" swimtime="00:01:31.56" />
                    <SPLIT distance="200" swimtime="00:01:45.67" />
                    <SPLIT distance="225" swimtime="00:01:58.28" />
                    <SPLIT distance="250" swimtime="00:02:12.30" />
                    <SPLIT distance="275" swimtime="00:02:26.43" />
                    <SPLIT distance="300" swimtime="00:02:40.23" />
                    <SPLIT distance="325" swimtime="00:02:52.07" />
                    <SPLIT distance="350" swimtime="00:03:05.61" />
                    <SPLIT distance="375" swimtime="00:03:19.55" />
                    <SPLIT distance="400" swimtime="00:03:33.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="165928" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="213597" reactiontime="+36" />
                    <RELAYPOSITION number="3" athleteid="202246" reactiontime="+36" />
                    <RELAYPOSITION number="4" athleteid="126805" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Great Britain">
              <RESULTS>
                <RESULT eventid="47" place="-1" lane="2" heat="1" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Great Britain">
              <RESULTS>
                <RESULT eventid="125" place="6" lane="2" heat="1" swimtime="00:01:37.11" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.57" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                    <SPLIT distance="75" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:00:48.31" />
                    <SPLIT distance="125" swimtime="00:00:59.70" />
                    <SPLIT distance="150" swimtime="00:01:12.49" />
                    <SPLIT distance="175" swimtime="00:01:24.18" />
                    <SPLIT distance="200" swimtime="00:01:37.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="165928" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="213597" reactiontime="+40" />
                    <RELAYPOSITION number="3" athleteid="161299" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="126805" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="5" lane="2" heat="2" swimtime="00:01:37.41" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:23.99" />
                    <SPLIT distance="75" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:00:48.18" />
                    <SPLIT distance="125" swimtime="00:00:59.86" />
                    <SPLIT distance="150" swimtime="00:01:12.78" />
                    <SPLIT distance="175" swimtime="00:01:24.49" />
                    <SPLIT distance="200" swimtime="00:01:37.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="165928" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="213597" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="161299" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="126805" reactiontime="+12" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Great Britain">
              <RESULTS>
                <RESULT eventid="34" place="-1" lane="8" heat="2" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Great Britain">
              <RESULTS>
                <RESULT eventid="111" place="4" lane="3" heat="1" swimtime="00:01:37.07" reactiontime="+80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                    <SPLIT distance="75" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:00:51.84" />
                    <SPLIT distance="125" swimtime="00:01:01.79" />
                    <SPLIT distance="150" swimtime="00:01:13.77" />
                    <SPLIT distance="175" swimtime="00:01:24.90" />
                    <SPLIT distance="200" swimtime="00:01:37.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202246" reactiontime="+80" />
                    <RELAYPOSITION number="2" athleteid="108588" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="101625" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="165928" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="3" lane="1" heat="3" swimtime="00:01:38.46" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:26.97" />
                    <SPLIT distance="75" swimtime="00:00:38.29" />
                    <SPLIT distance="100" swimtime="00:00:52.46" />
                    <SPLIT distance="125" swimtime="00:01:02.59" />
                    <SPLIT distance="150" swimtime="00:01:14.88" />
                    <SPLIT distance="175" swimtime="00:01:26.02" />
                    <SPLIT distance="200" swimtime="00:01:38.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202246" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="108588" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="101625" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="165928" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Georgia" shortname="GEO" code="GEO" nation="GEO" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198239" lastname="KUKHALASHVILI" firstname="Luka" gender="M" birthdate="2002-10-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.57" eventid="14" heat="6" lane="1">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:01:47.51" eventid="44" heat="2" lane="3">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="56" lane="1" heat="6" heatid="60014" swimtime="00:00:50.59" reactiontime="+66" points="696">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:24.12" />
                    <SPLIT distance="75" swimtime="00:00:37.37" />
                    <SPLIT distance="100" swimtime="00:00:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="37" lane="3" heat="2" heatid="20044" swimtime="00:01:49.38" reactiontime="+66" points="749">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:25.72" />
                    <SPLIT distance="75" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:00:53.40" />
                    <SPLIT distance="125" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:20.98" />
                    <SPLIT distance="175" swimtime="00:01:35.17" />
                    <SPLIT distance="200" swimtime="00:01:49.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197304" lastname="NIKOLAISHVILI" firstname="Salome" gender="F" birthdate="2006-03-26">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.97" eventid="2" heat="1" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.60" eventid="18" heat="3" lane="1">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="42" lane="4" heat="1" heatid="10002" swimtime="00:01:07.03" reactiontime="+55" points="549">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="75" swimtime="00:00:49.17" />
                    <SPLIT distance="100" swimtime="00:01:07.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="40" lane="1" heat="3" heatid="30018" swimtime="00:00:30.11" reactiontime="+55" points="591">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Germany" shortname="GER" code="GER" nation="GER" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="125264" lastname="ULRICH" firstname="Marek" gender="M" birthdate="1997-01-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.54" eventid="3" heat="3" lane="7">
                  <MEETINFO date="2021-07-26" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.49" eventid="19" heat="4" lane="2">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="16" lane="7" heat="3" heatid="30003" swimtime="00:00:50.92" reactiontime="+67" points="855">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:24.68" />
                    <SPLIT distance="75" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:00:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="16" lane="8" heat="1" heatid="10203" swimtime="00:00:51.12" reactiontime="+65" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.79" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:00:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="8" lane="1" heat="1" heatid="10119" swimtime="00:00:23.37" reactiontime="+65" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="14" lane="2" heat="4" heatid="40019" swimtime="00:00:23.28" reactiontime="+62" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="7" lane="1" heat="1" heatid="10219" swimtime="00:00:23.03" reactiontime="+59" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:23.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195394" lastname="BRAUNSCHWEIG" firstname="Ole" gender="M" birthdate="1997-11-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.69" eventid="3" heat="4" lane="6">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.28" eventid="19" heat="4" lane="6">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="10" lane="6" heat="4" heatid="40003" swimtime="00:00:50.37" reactiontime="+56" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="75" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:00:50.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="12" lane="2" heat="1" heatid="10203" swimtime="00:00:50.55" reactiontime="+60" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:24.35" />
                    <SPLIT distance="75" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:00:50.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="11" lane="6" heat="4" heatid="40019" swimtime="00:00:23.25" reactiontime="+57" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.47" />
                    <SPLIT distance="50" swimtime="00:00:23.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="11" lane="7" heat="2" heatid="20219" swimtime="00:00:23.08" reactiontime="+55" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.34" />
                    <SPLIT distance="50" swimtime="00:00:23.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195395" lastname="MATZERATH" firstname="Lucas" gender="M" birthdate="2000-05-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.57" eventid="16" heat="7" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:26.50" eventid="41" heat="9" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="7" lane="1" heat="1" heatid="10116" swimtime="00:00:57.12" reactiontime="+67" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:00:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="8" lane="1" heat="7" heatid="70016" swimtime="00:00:57.22" reactiontime="+68" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="75" swimtime="00:00:41.88" />
                    <SPLIT distance="100" swimtime="00:00:57.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="7" lane="6" heat="1" heatid="10216" swimtime="00:00:57.04" reactiontime="+66" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="75" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="19" lane="1" heat="9" heatid="90041" swimtime="00:00:26.67" reactiontime="+66" points="818">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="131055" lastname="KUSCH" firstname="Marius" gender="M" birthdate="1993-05-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.49" eventid="39" heat="8" lane="5">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.32" eventid="5" heat="10" lane="6">
                  <MEETINFO date="2021-09-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="3" lane="6" heat="1" heatid="10139" swimtime="00:00:49.12" reactiontime="+65" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:22.76" />
                    <SPLIT distance="75" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:00:49.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="7" lane="5" heat="8" heatid="80039" swimtime="00:00:49.89" reactiontime="+64" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.47" />
                    <SPLIT distance="50" swimtime="00:00:23.13" />
                    <SPLIT distance="75" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:00:49.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="4" lane="6" heat="2" heatid="20239" swimtime="00:00:49.20" reactiontime="+65" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.30" />
                    <SPLIT distance="50" swimtime="00:00:23.01" />
                    <SPLIT distance="75" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:00:49.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="105" place="7" lane="7" heat="1" heatid="10105" swimtime="00:00:22.17" reactiontime="+66" points="944">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.06" />
                    <SPLIT distance="50" swimtime="00:00:22.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="5" lane="6" heat="10" heatid="100005" swimtime="00:00:22.19" reactiontime="+64" points="941">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.05" />
                    <SPLIT distance="50" swimtime="00:00:22.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="6" lane="3" heat="2" heatid="20205" swimtime="00:00:22.14" reactiontime="+66" points="948">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:22.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149729" lastname="SALCHOW" firstname="Josha" gender="M" birthdate="1999-07-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.87" eventid="14" heat="10" lane="7">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.06" eventid="44" heat="6" lane="8">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:21.91" eventid="31" heat="7" lane="5">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="19" lane="7" heat="10" heatid="100014" swimtime="00:00:47.11" reactiontime="+71" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.60" />
                    <SPLIT distance="50" swimtime="00:00:22.46" />
                    <SPLIT distance="75" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="24" lane="8" heat="6" heatid="60044" swimtime="00:01:45.01" reactiontime="+72" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:24.57" />
                    <SPLIT distance="75" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:00:51.11" />
                    <SPLIT distance="125" swimtime="00:01:04.62" />
                    <SPLIT distance="150" swimtime="00:01:18.23" />
                    <SPLIT distance="175" swimtime="00:01:31.82" />
                    <SPLIT distance="200" swimtime="00:01:45.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="31" lane="5" heat="7" heatid="70031" swimtime="00:00:21.52" reactiontime="+68" points="822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:21.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101365" lastname="KOCH" firstname="Marco" gender="M" birthdate="1990-01-25">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.36" eventid="29" heat="5" lane="6">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="129" place="7" lane="1" heat="1" heatid="10129" swimtime="00:02:05.01" reactiontime="+68" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.79" />
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="75" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:01:00.18" />
                    <SPLIT distance="125" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:01:32.20" />
                    <SPLIT distance="175" swimtime="00:01:48.60" />
                    <SPLIT distance="200" swimtime="00:02:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="7" lane="6" heat="5" heatid="50029" swimtime="00:02:04.08" reactiontime="+67" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="75" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:00.15" />
                    <SPLIT distance="125" swimtime="00:01:16.23" />
                    <SPLIT distance="150" swimtime="00:01:32.00" />
                    <SPLIT distance="175" swimtime="00:01:48.05" />
                    <SPLIT distance="200" swimtime="00:02:04.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164531" lastname="ELENDT" firstname="Anna" gender="F" birthdate="2001-09-04">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.07" eventid="15" heat="5" lane="5">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.33" eventid="28" heat="4" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.10" eventid="40" heat="6" lane="7">
                  <MEETINFO date="2022-05-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="3" lane="8" heat="1" heatid="10115" swimtime="00:01:04.05" reactiontime="+69" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="75" swimtime="00:00:46.68" />
                    <SPLIT distance="100" swimtime="00:01:04.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="6" lane="5" heat="5" heatid="50015" swimtime="00:01:04.53" reactiontime="+72" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.95" />
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="75" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:04.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="8" lane="3" heat="1" heatid="10215" swimtime="00:01:04.46" reactiontime="+71" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.17" />
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="75" swimtime="00:00:47.14" />
                    <SPLIT distance="100" swimtime="00:01:04.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="-1" lane="2" heat="4" heatid="40028" swimtime="NT" status="DNS" />
                <RESULT eventid="140" place="5" lane="1" heat="1" heatid="10140" swimtime="00:00:29.30" reactiontime="+67" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.36" />
                    <SPLIT distance="50" swimtime="00:00:29.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="6" lane="7" heat="6" heatid="60040" swimtime="00:00:29.59" reactiontime="+70" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="7" lane="3" heat="1" heatid="10240" swimtime="00:00:29.52" reactiontime="+68" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149821" lastname="KÖHLER" firstname="Angelina" gender="F" birthdate="2000-11-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.90" eventid="38" heat="2" lane="7">
                  <MEETINFO date="2022-08-15" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.21" eventid="4" heat="6" lane="1">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="138" place="4" lane="6" heat="1" heatid="10138" swimtime="00:00:56.20" reactiontime="+71" points="916">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                    <SPLIT distance="75" swimtime="00:00:41.06" />
                    <SPLIT distance="100" swimtime="00:00:56.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="5" lane="7" heat="2" heatid="20038" swimtime="00:00:56.56" reactiontime="+74" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                    <SPLIT distance="75" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="4" lane="3" heat="2" heatid="20238" swimtime="00:00:56.23" reactiontime="+73" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                    <SPLIT distance="50" swimtime="00:00:26.29" />
                    <SPLIT distance="75" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:00:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="17" lane="1" heat="6" heatid="60004" swimtime="00:00:25.85" reactiontime="+70" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.95" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="304" place="19" lane="5" heat="1" heatid="10304" swimtime="00:00:26.05" reactiontime="+71" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Germany">
              <RESULTS>
                <RESULT eventid="148" place="5" lane="6" heat="1" swimtime="00:03:23.04" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                    <SPLIT distance="50" swimtime="00:00:24.25" />
                    <SPLIT distance="75" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:00:50.68" />
                    <SPLIT distance="125" swimtime="00:01:02.54" />
                    <SPLIT distance="150" swimtime="00:01:16.88" />
                    <SPLIT distance="175" swimtime="00:01:31.98" />
                    <SPLIT distance="200" swimtime="00:01:47.64" />
                    <SPLIT distance="225" swimtime="00:01:57.60" />
                    <SPLIT distance="250" swimtime="00:02:10.26" />
                    <SPLIT distance="275" swimtime="00:02:22.95" />
                    <SPLIT distance="300" swimtime="00:02:36.36" />
                    <SPLIT distance="325" swimtime="00:02:46.52" />
                    <SPLIT distance="350" swimtime="00:02:58.42" />
                    <SPLIT distance="375" swimtime="00:03:10.81" />
                    <SPLIT distance="400" swimtime="00:03:23.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="195394" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="195395" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="131055" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="149729" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="4" lane="7" heat="2" swimtime="00:03:24.51" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:24.42" />
                    <SPLIT distance="75" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:00:50.63" />
                    <SPLIT distance="125" swimtime="00:01:02.79" />
                    <SPLIT distance="150" swimtime="00:01:17.65" />
                    <SPLIT distance="175" swimtime="00:01:32.91" />
                    <SPLIT distance="200" swimtime="00:01:48.40" />
                    <SPLIT distance="225" swimtime="00:01:58.44" />
                    <SPLIT distance="250" swimtime="00:02:11.10" />
                    <SPLIT distance="275" swimtime="00:02:24.22" />
                    <SPLIT distance="300" swimtime="00:02:37.84" />
                    <SPLIT distance="325" swimtime="00:02:48.03" />
                    <SPLIT distance="350" swimtime="00:02:59.88" />
                    <SPLIT distance="375" swimtime="00:03:12.13" />
                    <SPLIT distance="400" swimtime="00:03:24.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="195394" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="195395" reactiontime="+41" />
                    <RELAYPOSITION number="3" athleteid="131055" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="149729" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Germany">
              <RESULTS>
                <RESULT eventid="111" place="-1" lane="5" heat="1" status="DSQ" swimtime="00:01:36.61" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:22.98" />
                    <SPLIT distance="75" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:00:51.65" />
                    <SPLIT distance="125" swimtime="00:01:01.11" />
                    <SPLIT distance="150" swimtime="00:01:13.15" />
                    <SPLIT distance="175" swimtime="00:01:24.22" />
                    <SPLIT distance="200" swimtime="00:01:36.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="195394" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="164531" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="131055" reactiontime="-6" status="DSQ" />
                    <RELAYPOSITION number="4" athleteid="149821" reactiontime="+17" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="2" lane="5" heat="3" swimtime="00:01:37.90" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:23.29" />
                    <SPLIT distance="75" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                    <SPLIT distance="125" swimtime="00:01:02.11" />
                    <SPLIT distance="150" swimtime="00:01:14.10" />
                    <SPLIT distance="175" swimtime="00:01:25.37" />
                    <SPLIT distance="200" swimtime="00:01:37.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="195394" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="164531" reactiontime="+27" />
                    <RELAYPOSITION number="3" athleteid="131055" reactiontime="-1" />
                    <RELAYPOSITION number="4" athleteid="149821" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Germany">
              <RESULTS>
                <RESULT eventid="135" place="6" lane="3" heat="1" swimtime="00:01:31.79" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:23.09" />
                    <SPLIT distance="75" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:00:48.96" />
                    <SPLIT distance="125" swimtime="00:00:58.69" />
                    <SPLIT distance="150" swimtime="00:01:10.68" />
                    <SPLIT distance="175" swimtime="00:01:20.56" />
                    <SPLIT distance="200" swimtime="00:01:31.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="195394" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="195395" reactiontime="+44" />
                    <RELAYPOSITION number="3" athleteid="131055" reactiontime="+21" />
                    <RELAYPOSITION number="4" athleteid="149729" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="3" lane="1" heat="3" swimtime="00:01:32.56" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:23.26" />
                    <SPLIT distance="75" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:00:49.41" />
                    <SPLIT distance="125" swimtime="00:00:59.38" />
                    <SPLIT distance="150" swimtime="00:01:11.41" />
                    <SPLIT distance="175" swimtime="00:01:21.30" />
                    <SPLIT distance="200" swimtime="00:01:32.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="125264" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="195395" reactiontime="+39" />
                    <RELAYPOSITION number="3" athleteid="131055" reactiontime="+33" />
                    <RELAYPOSITION number="4" athleteid="149729" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Ghana" shortname="GHA" code="GHA" nation="GHA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="106848" lastname="JACKSON" firstname="Abeku" gender="M" birthdate="2000-04-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.39" eventid="39" heat="4" lane="7">
                  <MEETINFO date="2021-07-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.08" eventid="5" heat="4" lane="4">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="34" lane="7" heat="4" heatid="40039" swimtime="00:00:52.36" reactiontime="+63" points="759">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.24" />
                    <SPLIT distance="50" swimtime="00:00:24.61" />
                    <SPLIT distance="75" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="50" lane="4" heat="4" heatid="40005" swimtime="00:00:23.87" reactiontime="+64" points="756">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.92" />
                    <SPLIT distance="50" swimtime="00:00:23.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197900" lastname="ADJEI" firstname="Nubia" gender="F" birthdate="2003-01-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.09" eventid="18" heat="3" lane="2">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.31" eventid="4" heat="2" lane="4">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="39" lane="2" heat="3" heatid="30018" swimtime="00:00:29.96" reactiontime="+59" points="600">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.85" />
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="33" lane="4" heat="2" heatid="20004" swimtime="00:00:29.11" reactiontime="+72" points="587">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.50" />
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Gibraltar" shortname="GIB" code="GIB" nation="GIB" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198025" lastname="CARROLL" firstname="Aidan" gender="M" birthdate="2000-07-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.17" eventid="39" heat="2" lane="4">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.84" eventid="5" heat="3" lane="4">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="45" lane="4" heat="2" heatid="20039" swimtime="00:00:56.02" reactiontime="+57" points="620">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:26.01" />
                    <SPLIT distance="75" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:00:56.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="-1" lane="4" heat="3" heatid="30005" swimtime="00:00:25.53" status="DSQ" reactiontime="+62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128923" lastname="SAVITZ" firstname="Matt Dylan" gender="M" birthdate="1999-01-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.53" eventid="14" heat="2" lane="5">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="00:01:58.69" eventid="44" heat="1" lane="6">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="69" lane="5" heat="2" heatid="20014" swimtime="00:00:53.37" reactiontime="+71" points="593">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.15" />
                    <SPLIT distance="50" swimtime="00:00:25.48" />
                    <SPLIT distance="75" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:00:53.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="42" lane="6" heat="1" heatid="10044" swimtime="00:01:54.02" reactiontime="+67" points="661">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="75" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:00:56.19" />
                    <SPLIT distance="125" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:25.47" />
                    <SPLIT distance="175" swimtime="00:01:40.01" />
                    <SPLIT distance="200" swimtime="00:01:54.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201463" lastname="KENT" firstname="Asia" gender="F" birthdate="2007-03-13">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.80" eventid="15" heat="2" lane="7">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:02:43.98" eventid="28" heat="1" lane="6">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="43" lane="7" heat="2" heatid="20015" swimtime="00:01:13.80" reactiontime="+72" points="603">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="75" swimtime="00:00:53.56" />
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="29" lane="6" heat="1" heatid="10028" swimtime="00:02:36.22" reactiontime="+68" points="639">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.92" />
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="75" swimtime="00:00:53.66" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="125" swimtime="00:01:34.12" />
                    <SPLIT distance="150" swimtime="00:01:54.54" />
                    <SPLIT distance="175" swimtime="00:02:15.46" />
                    <SPLIT distance="200" swimtime="00:02:36.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201461" lastname="SANDERS" firstname="Rachel" gender="F" birthdate="2004-12-06">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="4" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="38" lane="3" heat="1" heatid="10004" swimtime="00:00:31.29" reactiontime="+79" points="473">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.49" />
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="44" lane="5" heat="1" heatid="10030" swimtime="00:00:28.73" reactiontime="+76" points="508">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Greece" shortname="GRE" code="GRE" nation="GRE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="110744" lastname="CHRISTOU" firstname="Apostolos" gender="M" birthdate="1996-11-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.87" eventid="3" heat="6" lane="3">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.87" eventid="19" heat="6" lane="5">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="5" lane="6" heat="1" heatid="10103" swimtime="00:00:49.68" reactiontime="+59" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.54" />
                    <SPLIT distance="50" swimtime="00:00:23.83" />
                    <SPLIT distance="75" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:00:49.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="3" lane="3" heat="6" heatid="60003" swimtime="00:00:50.01" reactiontime="+56" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:23.69" />
                    <SPLIT distance="75" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="4" lane="5" heat="2" heatid="20203" swimtime="00:00:49.66" reactiontime="+57" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:23.92" />
                    <SPLIT distance="75" swimtime="00:00:36.88" />
                    <SPLIT distance="100" swimtime="00:00:49.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="6" lane="8" heat="1" heatid="10119" swimtime="00:00:23.10" reactiontime="+61" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.27" />
                    <SPLIT distance="50" swimtime="00:00:23.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="8" lane="5" heat="6" heatid="60019" swimtime="00:00:23.18" reactiontime="+57" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                    <SPLIT distance="50" swimtime="00:00:23.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="8" lane="6" heat="1" heatid="10219" swimtime="00:00:23.05" reactiontime="+58" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.33" />
                    <SPLIT distance="50" swimtime="00:00:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="419" place="8" lane="4" heat="1" heatid="10419" swimtime="00:00:23.15" reactiontime="+56" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:23.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110782" lastname="VAZAIOS" firstname="Andreas" gender="M" birthdate="1994-05-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.35" eventid="21" heat="4" lane="6">
                  <MEETINFO date="2021-09-05" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.15" eventid="7" heat="3" lane="4">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:04:03.37" eventid="37" heat="2" lane="6">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.54" eventid="23" heat="3" lane="5">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="21" place="12" lane="6" heat="4" heatid="40021" swimtime="00:01:52.28" reactiontime="+65" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:25.52" />
                    <SPLIT distance="75" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:00:54.23" />
                    <SPLIT distance="125" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:22.77" />
                    <SPLIT distance="175" swimtime="00:01:37.17" />
                    <SPLIT distance="200" swimtime="00:01:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="10" lane="4" heat="3" heatid="30007" swimtime="00:01:53.08" reactiontime="+59" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:24.85" />
                    <SPLIT distance="75" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:00:52.66" />
                    <SPLIT distance="125" swimtime="00:01:09.08" />
                    <SPLIT distance="150" swimtime="00:01:25.73" />
                    <SPLIT distance="175" swimtime="00:01:39.89" />
                    <SPLIT distance="200" swimtime="00:01:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="16" lane="6" heat="2" heatid="20037" swimtime="00:04:11.39" reactiontime="+64" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                    <SPLIT distance="75" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                    <SPLIT distance="125" swimtime="00:01:12.40" />
                    <SPLIT distance="150" swimtime="00:01:27.94" />
                    <SPLIT distance="175" swimtime="00:01:43.73" />
                    <SPLIT distance="200" swimtime="00:01:59.04" />
                    <SPLIT distance="225" swimtime="00:02:16.20" />
                    <SPLIT distance="250" swimtime="00:02:33.45" />
                    <SPLIT distance="275" swimtime="00:02:51.22" />
                    <SPLIT distance="300" swimtime="00:03:09.37" />
                    <SPLIT distance="325" swimtime="00:03:24.90" />
                    <SPLIT distance="350" swimtime="00:03:40.42" />
                    <SPLIT distance="375" swimtime="00:03:56.18" />
                    <SPLIT distance="400" swimtime="00:04:11.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="6" lane="6" heat="1" heatid="10123" swimtime="00:00:51.80" reactiontime="+63" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.69" />
                    <SPLIT distance="50" swimtime="00:00:23.54" />
                    <SPLIT distance="75" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:00:51.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="14" lane="5" heat="3" heatid="30023" swimtime="00:00:52.62" reactiontime="+61" points="821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.94" />
                    <SPLIT distance="50" swimtime="00:00:24.03" />
                    <SPLIT distance="75" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:00:52.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="4" lane="1" heat="1" heatid="10223" swimtime="00:00:51.47" reactiontime="+62" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.39" />
                    <SPLIT distance="75" swimtime="00:00:38.60" />
                    <SPLIT distance="100" swimtime="00:00:51.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100976" lastname="GKOLOMEEV" firstname="Kristian" gender="M" birthdate="1993-07-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.14" eventid="5" heat="7" lane="7">
                  <MEETINFO date="2021-12-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.00" eventid="31" heat="9" lane="5">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="38" lane="7" heat="7" heatid="70005" swimtime="00:00:23.30" reactiontime="+68" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.55" />
                    <SPLIT distance="50" swimtime="00:00:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="14" lane="5" heat="9" heatid="90031" swimtime="00:00:21.21" reactiontime="+67" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.25" />
                    <SPLIT distance="50" swimtime="00:00:21.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="10" lane="1" heat="2" heatid="20231" swimtime="00:00:21.08" reactiontime="+66" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.15" />
                    <SPLIT distance="50" swimtime="00:00:21.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Guatemala" shortname="GUA" code="GUA" nation="GUA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="213802" lastname="VÁSQUEZ" firstname="Miguel" gender="M" birthdate="2000-08-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.45" eventid="14" heat="4" lane="1">
                  <MEETINFO date="2022-04-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.65" eventid="19" heat="1" lane="3">
                  <MEETINFO date="2022-04-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="50" lane="1" heat="4" heatid="40014" swimtime="00:00:49.77" reactiontime="+65" points="731">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:23.87" />
                    <SPLIT distance="75" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:00:49.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="35" lane="3" heat="1" heatid="10019" swimtime="00:00:25.31" reactiontime="+60" points="676">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:25.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155015" lastname="GORDILLO" firstname="Erick" gender="M" birthdate="1999-10-05">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.35" eventid="21" heat="3" lane="8">
                  <MEETINFO date="2022-04-24" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.47" eventid="7" heat="2" lane="7">
                  <MEETINFO date="2021-11-29" />
                </ENTRY>
                <ENTRY entrytime="00:04:14.58" eventid="37" heat="1" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="21" place="21" lane="8" heat="3" heatid="30021" swimtime="00:01:56.93" reactiontime="+63" points="793">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:55.16" />
                    <SPLIT distance="125" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:25.29" />
                    <SPLIT distance="175" swimtime="00:01:41.13" />
                    <SPLIT distance="200" swimtime="00:01:56.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="27" lane="7" heat="2" heatid="20007" swimtime="00:01:58.98" reactiontime="+64" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:25.41" />
                    <SPLIT distance="75" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:00:54.97" />
                    <SPLIT distance="125" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:29.88" />
                    <SPLIT distance="175" swimtime="00:01:44.95" />
                    <SPLIT distance="200" swimtime="00:01:58.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="15" lane="5" heat="1" heatid="10037" swimtime="00:04:10.97" reactiontime="+68" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:00:57.89" />
                    <SPLIT distance="125" swimtime="00:01:14.12" />
                    <SPLIT distance="150" swimtime="00:01:29.68" />
                    <SPLIT distance="175" swimtime="00:01:45.39" />
                    <SPLIT distance="200" swimtime="00:02:00.87" />
                    <SPLIT distance="225" swimtime="00:02:18.76" />
                    <SPLIT distance="250" swimtime="00:02:36.32" />
                    <SPLIT distance="275" swimtime="00:02:54.33" />
                    <SPLIT distance="300" swimtime="00:03:12.59" />
                    <SPLIT distance="325" swimtime="00:03:27.65" />
                    <SPLIT distance="350" swimtime="00:03:42.15" />
                    <SPLIT distance="375" swimtime="00:03:56.76" />
                    <SPLIT distance="400" swimtime="00:04:10.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="172253" lastname="JURADO" firstname="Krista" gender="F" birthdate="2004-01-06">
              <ENTRIES>
                <ENTRY entrytime="00:01:12.51" eventid="15" heat="3" lane="8">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:36.40" eventid="28" heat="1" lane="3">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="46" lane="8" heat="3" heatid="30015" swimtime="00:01:14.13" reactiontime="+70" points="595">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="75" swimtime="00:00:54.15" />
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="30" lane="3" heat="1" heatid="10028" swimtime="00:02:36.34" reactiontime="+66" points="637">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="75" swimtime="00:00:54.10" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="125" swimtime="00:01:34.35" />
                    <SPLIT distance="150" swimtime="00:01:54.93" />
                    <SPLIT distance="175" swimtime="00:02:15.55" />
                    <SPLIT distance="200" swimtime="00:02:36.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202424" lastname="MEJIA" firstname="Lucero" gender="F" birthdate="2007-10-17">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.78" eventid="43" heat="2" lane="8">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="00:05:03.61" eventid="36" heat="1" lane="5">
                  <MEETINFO date="2022-04-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="26" lane="8" heat="2" heatid="20043" swimtime="00:02:02.57" reactiontime="+66" points="728">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.36" />
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                    <SPLIT distance="75" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:00:59.88" />
                    <SPLIT distance="125" swimtime="00:01:15.74" />
                    <SPLIT distance="150" swimtime="00:01:31.52" />
                    <SPLIT distance="175" swimtime="00:01:47.34" />
                    <SPLIT distance="200" swimtime="00:02:02.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="22" lane="5" heat="1" heatid="10036" swimtime="00:04:49.99" reactiontime="+64" points="711">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="75" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                    <SPLIT distance="125" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:01:41.09" />
                    <SPLIT distance="175" swimtime="00:01:59.00" />
                    <SPLIT distance="200" swimtime="00:02:16.14" />
                    <SPLIT distance="225" swimtime="00:02:38.14" />
                    <SPLIT distance="250" swimtime="00:02:59.99" />
                    <SPLIT distance="275" swimtime="00:03:21.65" />
                    <SPLIT distance="300" swimtime="00:03:43.30" />
                    <SPLIT distance="325" swimtime="00:04:00.40" />
                    <SPLIT distance="350" swimtime="00:04:17.20" />
                    <SPLIT distance="375" swimtime="00:04:34.15" />
                    <SPLIT distance="400" swimtime="00:04:49.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Guatemala">
              <RESULTS>
                <RESULT eventid="11" place="25" lane="7" heat="1" swimtime="00:01:50.21" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.31" />
                    <SPLIT distance="50" swimtime="00:00:25.18" />
                    <SPLIT distance="75" swimtime="00:00:40.57" />
                    <SPLIT distance="100" swimtime="00:00:59.43" />
                    <SPLIT distance="125" swimtime="00:01:10.58" />
                    <SPLIT distance="150" swimtime="00:01:24.10" />
                    <SPLIT distance="175" swimtime="00:01:36.66" />
                    <SPLIT distance="200" swimtime="00:01:50.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213802" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="172253" reactiontime="+61" />
                    <RELAYPOSITION number="3" athleteid="155015" reactiontime="+49" />
                    <RELAYPOSITION number="4" athleteid="202424" reactiontime="+49" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Guinea" shortname="GUI" code="GUI" nation="GUI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197224" lastname="DIALLO" firstname="Elhadj N'gnane" gender="M" birthdate="2003-06-15">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.30" eventid="39" heat="2" lane="7">
                  <MEETINFO date="2022-08-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="55" lane="7" heat="2" heatid="20039" swimtime="00:01:05.58" reactiontime="+67" points="386">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                    <SPLIT distance="75" swimtime="00:00:46.77" />
                    <SPLIT distance="100" swimtime="00:01:05.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197220" lastname="CAMARA" firstname="Fode Amara" gender="M" birthdate="2005-01-01">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="14" heat="1" lane="7" />
                <ENTRY entrytime="00:00:27.84" eventid="31" heat="2" lane="4">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="-1" lane="7" heat="1" heatid="10014" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="-1" lane="4" heat="2" heatid="20031" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130109" lastname="TOURE" firstname="Mariama" gender="F" birthdate="2003-11-10">
              <ENTRIES>
                <ENTRY entrytime="00:01:36.59" eventid="15" heat="1" lane="5" />
                <ENTRY entrytime="00:00:41.91" eventid="40" heat="2" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="50" lane="5" heat="1" heatid="10015" swimtime="00:01:33.89" reactiontime="+70" points="292">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.10" />
                    <SPLIT distance="50" swimtime="00:00:42.19" />
                    <SPLIT distance="75" swimtime="00:01:07.63" />
                    <SPLIT distance="100" swimtime="00:01:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="40" lane="6" heat="2" heatid="20040" swimtime="00:00:40.92" reactiontime="+70" points="339">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.14" />
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Guam" shortname="GUM" code="GUM" nation="GUM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="159169" lastname="HENDRIX" firstname="James" gender="M" birthdate="2002-06-10">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="39" heat="2" lane="8" />
                <ENTRY entrytime="NT" eventid="21" heat="1" lane="6" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="46" lane="8" heat="2" heatid="20039" swimtime="00:00:56.08" reactiontime="+69" points="618">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:25.56" />
                    <SPLIT distance="75" swimtime="00:00:40.29" />
                    <SPLIT distance="100" swimtime="00:00:56.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="26" lane="6" heat="1" heatid="10021" swimtime="00:02:08.63" reactiontime="+72" points="595">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.23" />
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="75" swimtime="00:00:45.34" />
                    <SPLIT distance="100" swimtime="00:01:01.83" />
                    <SPLIT distance="125" swimtime="00:01:18.41" />
                    <SPLIT distance="150" swimtime="00:01:35.24" />
                    <SPLIT distance="175" swimtime="00:01:51.95" />
                    <SPLIT distance="200" swimtime="00:02:08.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197804" lastname="POPPE" firstname="Israel" gender="M" birthdate="2006-11-26">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.89" eventid="44" heat="1" lane="2">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="24" heat="1" lane="1" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="44" lane="2" heat="1" heatid="10044" swimtime="00:01:57.67" reactiontime="+59" points="602">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.44" />
                    <SPLIT distance="50" swimtime="00:00:26.75" />
                    <SPLIT distance="75" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:00:57.13" />
                    <SPLIT distance="125" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:27.52" />
                    <SPLIT distance="175" swimtime="00:01:43.00" />
                    <SPLIT distance="200" swimtime="00:01:57.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="34" lane="1" heat="1" heatid="10024" swimtime="00:04:17.65" reactiontime="+61" points="559">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                    <SPLIT distance="75" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:00:59.39" />
                    <SPLIT distance="125" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:31.63" />
                    <SPLIT distance="175" swimtime="00:01:48.04" />
                    <SPLIT distance="200" swimtime="00:02:04.33" />
                    <SPLIT distance="225" swimtime="00:02:20.79" />
                    <SPLIT distance="250" swimtime="00:02:37.41" />
                    <SPLIT distance="275" swimtime="00:02:54.04" />
                    <SPLIT distance="300" swimtime="00:03:10.91" />
                    <SPLIT distance="325" swimtime="00:03:27.90" />
                    <SPLIT distance="350" swimtime="00:03:44.93" />
                    <SPLIT distance="375" swimtime="00:04:01.81" />
                    <SPLIT distance="400" swimtime="00:04:17.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202092" lastname="LEE" firstname="Mia" gender="F" birthdate="2008-05-12">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:03.67" eventid="13" heat="2" lane="4">
                  <MEETINFO date="2022-06-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="52" lane="4" heat="2" heatid="20013" swimtime="00:01:00.38" reactiontime="+62" points="576">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="75" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="27" lane="3" heat="1" heatid="10022" swimtime="00:01:10.55" reactiontime="+66" points="513">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.19" />
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="75" swimtime="00:00:54.10" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214624" lastname="BOLLINGER" firstname="Amaya" gender="F" birthdate="2008-07-03">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="20" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="1" heat="1" lane="7" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="24" lane="3" heat="1" heatid="10020" swimtime="00:02:35.87" reactiontime="+76" points="451">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="75" swimtime="00:00:51.85" />
                    <SPLIT distance="100" swimtime="00:01:10.47" />
                    <SPLIT distance="125" swimtime="00:01:30.15" />
                    <SPLIT distance="150" swimtime="00:01:51.14" />
                    <SPLIT distance="175" swimtime="00:02:12.79" />
                    <SPLIT distance="200" swimtime="00:02:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="28" lane="7" heat="1" heatid="10001" swimtime="00:05:04.88" reactiontime="+70" points="451">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.52" />
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="75" swimtime="00:00:50.72" />
                    <SPLIT distance="100" swimtime="00:01:08.96" />
                    <SPLIT distance="125" swimtime="00:01:27.72" />
                    <SPLIT distance="150" swimtime="00:01:46.58" />
                    <SPLIT distance="175" swimtime="00:02:05.94" />
                    <SPLIT distance="200" swimtime="00:02:25.36" />
                    <SPLIT distance="225" swimtime="00:02:45.15" />
                    <SPLIT distance="250" swimtime="00:03:04.94" />
                    <SPLIT distance="275" swimtime="00:03:25.36" />
                    <SPLIT distance="300" swimtime="00:03:45.72" />
                    <SPLIT distance="325" swimtime="00:04:06.10" />
                    <SPLIT distance="350" swimtime="00:04:26.22" />
                    <SPLIT distance="375" swimtime="00:04:45.89" />
                    <SPLIT distance="400" swimtime="00:05:04.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Guam">
              <RESULTS>
                <RESULT eventid="27" place="21" lane="2" heat="3" swimtime="00:01:43.86" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:24.10" />
                    <SPLIT distance="75" swimtime="00:00:36.81" />
                    <SPLIT distance="100" swimtime="00:00:51.22" />
                    <SPLIT distance="125" swimtime="00:01:04.97" />
                    <SPLIT distance="150" swimtime="00:01:20.19" />
                    <SPLIT distance="175" swimtime="00:01:31.53" />
                    <SPLIT distance="200" swimtime="00:01:43.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="159169" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="202092" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="214624" reactiontime="+6" />
                    <RELAYPOSITION number="4" athleteid="197804" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Guam">
              <RESULTS>
                <RESULT eventid="11" place="30" lane="2" heat="1" swimtime="00:02:02.96" reactiontime="+82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.01" />
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="75" swimtime="00:00:52.96" />
                    <SPLIT distance="100" swimtime="00:01:13.28" />
                    <SPLIT distance="125" swimtime="00:01:25.27" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                    <SPLIT distance="175" swimtime="00:01:50.65" />
                    <SPLIT distance="200" swimtime="00:02:02.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214624" reactiontime="+82" />
                    <RELAYPOSITION number="2" athleteid="202092" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="159169" reactiontime="+46" />
                    <RELAYPOSITION number="4" athleteid="197804" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Guyana" shortname="GUY" code="GUY" nation="GUY" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="164034" lastname="SEATON" firstname="Leon" gender="M" birthdate="2004-05-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.56" eventid="14" heat="4" lane="4">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.85" eventid="31" heat="5" lane="8">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="61" lane="4" heat="4" heatid="40014" swimtime="00:00:51.24" reactiontime="+61" points="670">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:24.68" />
                    <SPLIT distance="75" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:00:51.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="54" lane="8" heat="5" heatid="50031" swimtime="00:00:23.65" reactiontime="+63" points="619">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.47" />
                    <SPLIT distance="50" swimtime="00:00:23.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197988" lastname="PERSAUD" firstname="Aleka Kylela" gender="F" birthdate="2006-02-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.70" eventid="13" heat="4" lane="1">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.86" eventid="30" heat="4" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="48" lane="1" heat="4" heatid="40013" swimtime="00:00:59.06" reactiontime="+57" points="615">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.02" />
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="75" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="36" lane="1" heat="4" heatid="40030" swimtime="00:00:26.42" reactiontime="+59" points="653">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Haiti" shortname="HAI" code="HAI" nation="HAI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="162310" lastname="GRAND'PIERRE" firstname="Alexandre" gender="M" birthdate="2003-01-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.34" eventid="16" heat="3" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.70" eventid="41" heat="3" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="47" lane="2" heat="3" heatid="30016" swimtime="00:01:01.07" reactiontime="+65" points="741">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="75" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:01.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="44" lane="4" heat="3" heatid="30041" swimtime="00:00:27.99" reactiontime="+64" points="708">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="160970" lastname="GRAND'PIERRE" firstname="Emilie Faith" gender="F" birthdate="2001-05-03">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.13" eventid="15" heat="2" lane="3">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.20" eventid="40" heat="3" lane="1">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="48" lane="3" heat="2" heatid="20015" swimtime="00:01:15.19" reactiontime="+68" points="570">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                    <SPLIT distance="75" swimtime="00:00:54.69" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="33" lane="1" heat="3" heatid="30040" swimtime="00:00:33.71" reactiontime="+68" points="608">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Hong Kong, China" shortname="HKG" code="HKG" nation="HKG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="151685" lastname="NG" firstname="Cheuk Yin" gender="M" birthdate="2002-09-25">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.87" eventid="3" heat="4" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.45" eventid="39" heat="5" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.68" eventid="19" heat="4" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.17" eventid="5" heat="7" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="20" lane="1" heat="4" heatid="40003" swimtime="00:00:51.30" reactiontime="+50" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                    <SPLIT distance="50" swimtime="00:00:24.42" />
                    <SPLIT distance="75" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:00:51.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="31" lane="1" heat="5" heatid="50039" swimtime="00:00:51.94" reactiontime="+66" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.96" />
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="75" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:00:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="25" lane="1" heat="4" heatid="40019" swimtime="00:00:23.83" reactiontime="+50" points="810">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:23.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="36" lane="1" heat="7" heatid="70005" swimtime="00:00:23.19" reactiontime="+64" points="825">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.78" />
                    <SPLIT distance="50" swimtime="00:00:23.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201488" lastname="CHILLINGWORTH" firstname="Adam John" gender="M" birthdate="1997-09-23">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.87" eventid="16" heat="4" lane="8">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.13" eventid="29" heat="4" lane="1">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="36" lane="8" heat="4" heatid="40016" swimtime="00:00:59.61" reactiontime="+67" points="797">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                    <SPLIT distance="75" swimtime="00:00:43.72" />
                    <SPLIT distance="100" swimtime="00:00:59.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="14" lane="1" heat="4" heatid="40029" swimtime="00:02:06.46" reactiontime="+63" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="75" swimtime="00:00:44.73" />
                    <SPLIT distance="100" swimtime="00:01:00.85" />
                    <SPLIT distance="125" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:01:33.49" />
                    <SPLIT distance="175" swimtime="00:01:50.11" />
                    <SPLIT distance="200" swimtime="00:02:06.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165123" lastname="HO" firstname="Ian Yentou" gender="M" birthdate="1997-04-25">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.08" eventid="14" heat="8" lane="1">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.22" eventid="31" heat="9" lane="2">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="33" lane="1" heat="8" heatid="80014" swimtime="00:00:47.61" reactiontime="+60" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.95" />
                    <SPLIT distance="50" swimtime="00:00:23.01" />
                    <SPLIT distance="75" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:00:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="5" lane="2" heat="9" heatid="90031" swimtime="00:00:20.99" reactiontime="+58" points="886">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.19" />
                    <SPLIT distance="50" swimtime="00:00:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="9" lane="3" heat="2" heatid="20231" swimtime="00:00:21.04" reactiontime="+59" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.20" />
                    <SPLIT distance="50" swimtime="00:00:21.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213133" lastname="KWAN" firstname="Hayden" gender="M" birthdate="2002-11-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:55.07" eventid="46" heat="2" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.70" eventid="7" heat="2" lane="2">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="18" lane="1" heat="2" heatid="20046" swimtime="00:01:53.95" reactiontime="+59" points="796">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:00:56.01" />
                    <SPLIT distance="125" swimtime="00:01:10.53" />
                    <SPLIT distance="150" swimtime="00:01:25.12" />
                    <SPLIT distance="175" swimtime="00:01:39.64" />
                    <SPLIT distance="200" swimtime="00:01:53.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="32" lane="2" heat="2" heatid="20007" swimtime="00:01:59.91" reactiontime="+68" points="764">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                    <SPLIT distance="75" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:00:54.47" />
                    <SPLIT distance="125" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:31.01" />
                    <SPLIT distance="175" swimtime="00:01:46.16" />
                    <SPLIT distance="200" swimtime="00:01:59.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129558" lastname="CHEUK" firstname="Ming Ho" gender="M" birthdate="2002-05-18">
              <ENTRIES>
                <ENTRY entrytime="00:01:46.50" eventid="44" heat="3" lane="7">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:03:47.51" eventid="24" heat="2" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="30" lane="7" heat="3" heatid="30044" swimtime="00:01:47.30" reactiontime="+63" points="794">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="75" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:00:52.62" />
                    <SPLIT distance="125" swimtime="00:01:06.35" />
                    <SPLIT distance="150" swimtime="00:01:20.21" />
                    <SPLIT distance="175" swimtime="00:01:33.89" />
                    <SPLIT distance="200" swimtime="00:01:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="25" lane="4" heat="2" heatid="20024" swimtime="00:03:49.94" reactiontime="+66" points="786">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.09" />
                    <SPLIT distance="50" swimtime="00:00:25.76" />
                    <SPLIT distance="75" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:00:54.13" />
                    <SPLIT distance="125" swimtime="00:01:08.29" />
                    <SPLIT distance="150" swimtime="00:01:22.74" />
                    <SPLIT distance="175" swimtime="00:01:37.24" />
                    <SPLIT distance="200" swimtime="00:01:51.73" />
                    <SPLIT distance="225" swimtime="00:02:06.45" />
                    <SPLIT distance="250" swimtime="00:02:21.29" />
                    <SPLIT distance="275" swimtime="00:02:36.21" />
                    <SPLIT distance="300" swimtime="00:02:51.23" />
                    <SPLIT distance="325" swimtime="00:03:06.18" />
                    <SPLIT distance="350" swimtime="00:03:21.04" />
                    <SPLIT distance="375" swimtime="00:03:35.90" />
                    <SPLIT distance="400" swimtime="00:03:49.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105413" lastname="NG" firstname="Yan Kin" gender="M" birthdate="1997-07-25">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:27.49" eventid="41" heat="5" lane="6">
                  <MEETINFO date="2021-09-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="43" lane="6" heat="5" heatid="50041" swimtime="00:00:27.92" reactiontime="+60" points="713">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101305" lastname="AU" firstname="Hoi Shun Stephanie" gender="F" birthdate="1992-05-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.79" eventid="2" heat="6" lane="8">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:27.42" eventid="18" heat="7" lane="8">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="28" lane="8" heat="6" heatid="60002" swimtime="00:00:59.05" reactiontime="+57" points="803">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.85" />
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                    <SPLIT distance="75" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:00:59.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="26" lane="8" heat="7" heatid="70018" swimtime="00:00:27.30" reactiontime="+59" points="793">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.45" />
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="151671" lastname="LAM" firstname="Hoi Kiu" gender="F" birthdate="2003-11-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:09.11" eventid="15" heat="3" lane="6">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:00:31.33" eventid="40" heat="4" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="36" lane="6" heat="3" heatid="30015" swimtime="00:01:09.04" reactiontime="+64" points="736">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.97" />
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="75" swimtime="00:00:50.55" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="28" lane="1" heat="4" heatid="40040" swimtime="00:00:31.71" reactiontime="+51" points="730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100989" lastname="SZE" firstname="Hang Yu" gender="F" birthdate="1988-03-05">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:59.03" eventid="38" heat="3" lane="8">
                  <MEETINFO date="2022-09-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="20" lane="8" heat="3" heatid="30038" swimtime="00:00:58.06" reactiontime="+70" points="831">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                    <SPLIT distance="75" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:00:58.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122606" lastname="HAUGHEY" firstname="Siobhan Bernadette" gender="F" birthdate="1997-10-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.79" eventid="13" heat="8" lane="4">
                  <MEETINFO date="2021-12-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.31" eventid="43" heat="5" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="2" lane="5" heat="1" heatid="10113" swimtime="00:00:50.87" reactiontime="+71" points="963">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:24.59" />
                    <SPLIT distance="75" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:00:50.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="1" lane="4" heat="8" heatid="80013" swimtime="00:00:52.04" reactiontime="+72" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:24.69" />
                    <SPLIT distance="75" swimtime="00:00:38.31" />
                    <SPLIT distance="100" swimtime="00:00:52.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="2" lane="4" heat="2" heatid="20213" swimtime="00:00:51.69" reactiontime="+76" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:25.08" />
                    <SPLIT distance="75" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="143" place="1" lane="5" heat="1" heatid="10143" swimtime="00:01:51.65" reactiontime="+71" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                    <SPLIT distance="75" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:00:54.30" />
                    <SPLIT distance="125" swimtime="00:01:08.54" />
                    <SPLIT distance="150" swimtime="00:01:22.79" />
                    <SPLIT distance="175" swimtime="00:01:37.16" />
                    <SPLIT distance="200" swimtime="00:01:51.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="2" lane="4" heat="5" heatid="50043" swimtime="00:01:53.39" reactiontime="+73" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                    <SPLIT distance="75" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:00:55.83" />
                    <SPLIT distance="125" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:24.66" />
                    <SPLIT distance="175" swimtime="00:01:39.18" />
                    <SPLIT distance="200" swimtime="00:01:53.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210408" lastname="CHEUNG" firstname="Sum Yuet Cindy" gender="F" birthdate="2006-08-09">
              <ENTRIES>
                <ENTRY entrytime="00:02:14.53" eventid="45" heat="2" lane="8">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="28" lane="8" heat="2" heatid="20045" swimtime="00:02:09.55" reactiontime="+60" points="773">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="75" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                    <SPLIT distance="125" swimtime="00:01:19.48" />
                    <SPLIT distance="150" swimtime="00:01:36.50" />
                    <SPLIT distance="175" swimtime="00:01:53.34" />
                    <SPLIT distance="200" swimtime="00:02:09.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214616" lastname="CHANG" firstname="Yujuan" gender="F" birthdate="2000-04-09">
              <ENTRIES>
                <ENTRY entrytime="00:02:27.45" eventid="28" heat="2" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="25" lane="1" heat="2" heatid="20028" swimtime="00:02:26.76" reactiontime="+71" points="770">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.43" />
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="75" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                    <SPLIT distance="125" swimtime="00:01:29.66" />
                    <SPLIT distance="150" swimtime="00:01:48.45" />
                    <SPLIT distance="175" swimtime="00:02:07.30" />
                    <SPLIT distance="200" swimtime="00:02:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="23" lane="7" heat="1" heatid="10022" swimtime="00:01:02.64" reactiontime="+74" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="75" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:02.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214617" lastname="YEUNG" firstname="Hoi Ching" gender="F" birthdate="2007-03-18">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.98" eventid="20" heat="4" lane="8">
                  <MEETINFO date="2022-09-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.71" eventid="6" heat="1" lane="4">
                  <MEETINFO date="2021-09-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="22" lane="8" heat="4" heatid="40020" swimtime="00:02:12.57" reactiontime="+71" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.26" />
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="75" swimtime="00:00:45.79" />
                    <SPLIT distance="100" swimtime="00:01:03.18" />
                    <SPLIT distance="125" swimtime="00:01:20.50" />
                    <SPLIT distance="150" swimtime="00:01:38.11" />
                    <SPLIT distance="175" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="32" lane="4" heat="1" heatid="10006" swimtime="00:02:19.41" reactiontime="+67" points="667">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="75" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                    <SPLIT distance="125" swimtime="00:01:25.97" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="175" swimtime="00:02:03.88" />
                    <SPLIT distance="200" swimtime="00:02:19.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129491" lastname="HO" firstname="Nam Wai Tinky" gender="F" birthdate="2002-04-30">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:04:13.10" eventid="1" heat="2" lane="1">
                  <MEETINFO date="2022-07-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="21" lane="1" heat="2" heatid="20001" swimtime="00:04:14.15" reactiontime="+71" points="779">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                    <SPLIT distance="75" swimtime="00:00:44.85" />
                    <SPLIT distance="100" swimtime="00:01:00.67" />
                    <SPLIT distance="125" swimtime="00:01:16.73" />
                    <SPLIT distance="150" swimtime="00:01:32.52" />
                    <SPLIT distance="175" swimtime="00:01:48.36" />
                    <SPLIT distance="200" swimtime="00:02:04.33" />
                    <SPLIT distance="225" swimtime="00:02:20.48" />
                    <SPLIT distance="250" swimtime="00:02:36.79" />
                    <SPLIT distance="275" swimtime="00:02:53.11" />
                    <SPLIT distance="300" swimtime="00:03:09.44" />
                    <SPLIT distance="325" swimtime="00:03:25.97" />
                    <SPLIT distance="350" swimtime="00:03:42.25" />
                    <SPLIT distance="375" swimtime="00:03:58.55" />
                    <SPLIT distance="400" swimtime="00:04:14.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210412" lastname="NG" firstname="Lai Wa" gender="F" birthdate="2005-10-08">
              <ENTRIES>
                <ENTRY entrytime="00:04:52.39" eventid="36" heat="1" lane="4">
                  <MEETINFO date="2021-08-08" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:17:21.71" eventid="33" heat="1" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="36" place="20" lane="4" heat="1" heatid="10036" swimtime="00:04:45.62" reactiontime="+54" points="745">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                    <SPLIT distance="75" swimtime="00:00:47.80" />
                    <SPLIT distance="100" swimtime="00:01:05.54" />
                    <SPLIT distance="125" swimtime="00:01:24.27" />
                    <SPLIT distance="150" swimtime="00:01:41.53" />
                    <SPLIT distance="175" swimtime="00:01:59.50" />
                    <SPLIT distance="200" swimtime="00:02:16.52" />
                    <SPLIT distance="225" swimtime="00:02:37.13" />
                    <SPLIT distance="250" swimtime="00:02:58.07" />
                    <SPLIT distance="275" swimtime="00:03:18.91" />
                    <SPLIT distance="300" swimtime="00:03:40.04" />
                    <SPLIT distance="325" swimtime="00:03:57.00" />
                    <SPLIT distance="350" swimtime="00:04:13.58" />
                    <SPLIT distance="375" swimtime="00:04:29.88" />
                    <SPLIT distance="400" swimtime="00:04:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="15" lane="3" heat="1" heatid="10033" swimtime="00:17:01.32" reactiontime="+66" points="726">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="75" swimtime="00:00:45.61" />
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="125" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:01:35.37" />
                    <SPLIT distance="175" swimtime="00:01:52.25" />
                    <SPLIT distance="200" swimtime="00:02:08.97" />
                    <SPLIT distance="225" swimtime="00:02:25.78" />
                    <SPLIT distance="250" swimtime="00:02:42.44" />
                    <SPLIT distance="275" swimtime="00:02:59.35" />
                    <SPLIT distance="300" swimtime="00:03:16.22" />
                    <SPLIT distance="325" swimtime="00:03:33.23" />
                    <SPLIT distance="350" swimtime="00:03:50.06" />
                    <SPLIT distance="375" swimtime="00:04:07.13" />
                    <SPLIT distance="400" swimtime="00:04:23.97" />
                    <SPLIT distance="425" swimtime="00:04:41.08" />
                    <SPLIT distance="450" swimtime="00:04:58.06" />
                    <SPLIT distance="475" swimtime="00:05:14.77" />
                    <SPLIT distance="500" swimtime="00:05:32.07" />
                    <SPLIT distance="525" swimtime="00:05:48.75" />
                    <SPLIT distance="550" swimtime="00:06:06.10" />
                    <SPLIT distance="575" swimtime="00:06:22.82" />
                    <SPLIT distance="600" swimtime="00:06:39.78" />
                    <SPLIT distance="625" swimtime="00:06:56.97" />
                    <SPLIT distance="650" swimtime="00:07:14.20" />
                    <SPLIT distance="675" swimtime="00:07:31.43" />
                    <SPLIT distance="700" swimtime="00:07:48.59" />
                    <SPLIT distance="725" swimtime="00:08:05.75" />
                    <SPLIT distance="750" swimtime="00:08:22.81" />
                    <SPLIT distance="775" swimtime="00:08:39.85" />
                    <SPLIT distance="800" swimtime="00:08:57.15" />
                    <SPLIT distance="825" swimtime="00:09:14.44" />
                    <SPLIT distance="850" swimtime="00:09:31.51" />
                    <SPLIT distance="875" swimtime="00:09:48.68" />
                    <SPLIT distance="900" swimtime="00:10:05.85" />
                    <SPLIT distance="925" swimtime="00:10:23.05" />
                    <SPLIT distance="950" swimtime="00:10:40.31" />
                    <SPLIT distance="975" swimtime="00:10:57.54" />
                    <SPLIT distance="1000" swimtime="00:11:15.01" />
                    <SPLIT distance="1025" swimtime="00:11:31.96" />
                    <SPLIT distance="1050" swimtime="00:11:49.43" />
                    <SPLIT distance="1075" swimtime="00:12:06.77" />
                    <SPLIT distance="1100" swimtime="00:12:24.11" />
                    <SPLIT distance="1125" swimtime="00:12:41.31" />
                    <SPLIT distance="1150" swimtime="00:12:58.69" />
                    <SPLIT distance="1175" swimtime="00:13:16.24" />
                    <SPLIT distance="1200" swimtime="00:13:33.54" />
                    <SPLIT distance="1225" swimtime="00:13:50.96" />
                    <SPLIT distance="1250" swimtime="00:14:08.26" />
                    <SPLIT distance="1275" swimtime="00:14:25.64" />
                    <SPLIT distance="1300" swimtime="00:14:42.92" />
                    <SPLIT distance="1325" swimtime="00:15:00.37" />
                    <SPLIT distance="1350" swimtime="00:15:17.80" />
                    <SPLIT distance="1375" swimtime="00:15:35.43" />
                    <SPLIT distance="1400" swimtime="00:15:53.09" />
                    <SPLIT distance="1425" swimtime="00:16:10.59" />
                    <SPLIT distance="1450" swimtime="00:16:27.71" />
                    <SPLIT distance="1475" swimtime="00:16:44.84" />
                    <SPLIT distance="1500" swimtime="00:17:01.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101068" lastname="CHAN" firstname="Kin Lok" gender="F" birthdate="1994-03-07">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:26.67" eventid="4" heat="4" lane="8">
                  <MEETINFO date="2021-09-12" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.31" eventid="30" heat="5" lane="3">
                  <MEETINFO date="2021-09-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="27" lane="8" heat="4" heatid="40004" swimtime="00:00:27.08" reactiontime="+69" points="729">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="30" lane="3" heat="5" heatid="50030" swimtime="00:00:25.61" reactiontime="+70" points="717">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                    <SPLIT distance="50" swimtime="00:00:25.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="9" place="11" lane="2" heat="1" swimtime="00:03:14.67" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.25" />
                    <SPLIT distance="50" swimtime="00:00:23.56" />
                    <SPLIT distance="75" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:00:48.71" />
                    <SPLIT distance="125" swimtime="00:00:59.28" />
                    <SPLIT distance="150" swimtime="00:01:11.24" />
                    <SPLIT distance="175" swimtime="00:01:23.80" />
                    <SPLIT distance="200" swimtime="00:01:36.66" />
                    <SPLIT distance="225" swimtime="00:01:47.67" />
                    <SPLIT distance="250" swimtime="00:02:00.36" />
                    <SPLIT distance="275" swimtime="00:02:13.54" />
                    <SPLIT distance="300" swimtime="00:02:26.83" />
                    <SPLIT distance="325" swimtime="00:02:37.04" />
                    <SPLIT distance="350" swimtime="00:02:49.31" />
                    <SPLIT distance="375" swimtime="00:03:01.98" />
                    <SPLIT distance="400" swimtime="00:03:14.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129558" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="165123" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="105413" reactiontime="+17" />
                    <RELAYPOSITION number="4" athleteid="151685" reactiontime="+4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="48" place="13" lane="8" heat="3" swimtime="00:03:30.73" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:00:52.96" />
                    <SPLIT distance="125" swimtime="00:01:05.73" />
                    <SPLIT distance="150" swimtime="00:01:20.89" />
                    <SPLIT distance="175" swimtime="00:01:36.46" />
                    <SPLIT distance="200" swimtime="00:01:52.37" />
                    <SPLIT distance="225" swimtime="00:02:02.84" />
                    <SPLIT distance="250" swimtime="00:02:15.62" />
                    <SPLIT distance="275" swimtime="00:02:29.11" />
                    <SPLIT distance="300" swimtime="00:02:43.50" />
                    <SPLIT distance="325" swimtime="00:02:53.57" />
                    <SPLIT distance="350" swimtime="00:03:05.62" />
                    <SPLIT distance="375" swimtime="00:03:18.06" />
                    <SPLIT distance="400" swimtime="00:03:30.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213133" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="201488" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="151685" reactiontime="+9" />
                    <RELAYPOSITION number="4" athleteid="165123" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="32" place="12" lane="7" heat="2" swimtime="00:07:21.61" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:24.72" />
                    <SPLIT distance="75" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:00:51.73" />
                    <SPLIT distance="125" swimtime="00:01:05.30" />
                    <SPLIT distance="150" swimtime="00:01:19.48" />
                    <SPLIT distance="175" swimtime="00:01:33.55" />
                    <SPLIT distance="200" swimtime="00:01:47.15" />
                    <SPLIT distance="225" swimtime="00:01:58.49" />
                    <SPLIT distance="250" swimtime="00:02:11.41" />
                    <SPLIT distance="275" swimtime="00:02:25.20" />
                    <SPLIT distance="300" swimtime="00:02:39.12" />
                    <SPLIT distance="325" swimtime="00:02:52.97" />
                    <SPLIT distance="350" swimtime="00:03:07.19" />
                    <SPLIT distance="375" swimtime="00:03:21.81" />
                    <SPLIT distance="400" swimtime="00:03:36.17" />
                    <SPLIT distance="425" swimtime="00:03:48.08" />
                    <SPLIT distance="450" swimtime="00:04:01.92" />
                    <SPLIT distance="475" swimtime="00:04:16.03" />
                    <SPLIT distance="500" swimtime="00:04:30.41" />
                    <SPLIT distance="525" swimtime="00:04:44.67" />
                    <SPLIT distance="550" swimtime="00:04:59.21" />
                    <SPLIT distance="575" swimtime="00:05:13.84" />
                    <SPLIT distance="600" swimtime="00:05:27.98" />
                    <SPLIT distance="625" swimtime="00:05:39.88" />
                    <SPLIT distance="650" swimtime="00:05:53.35" />
                    <SPLIT distance="675" swimtime="00:06:07.31" />
                    <SPLIT distance="700" swimtime="00:06:21.96" />
                    <SPLIT distance="725" swimtime="00:06:36.46" />
                    <SPLIT distance="750" swimtime="00:06:51.72" />
                    <SPLIT distance="775" swimtime="00:07:06.73" />
                    <SPLIT distance="800" swimtime="00:07:21.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129558" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="213133" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="201488" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="105413" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="26" place="11" lane="3" heat="1" swimtime="00:01:27.59" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.04" />
                    <SPLIT distance="50" swimtime="00:00:22.93" />
                    <SPLIT distance="75" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:00:43.88" />
                    <SPLIT distance="125" swimtime="00:00:53.95" />
                    <SPLIT distance="150" swimtime="00:01:05.24" />
                    <SPLIT distance="175" swimtime="00:01:16.08" />
                    <SPLIT distance="200" swimtime="00:01:27.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129558" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="165123" reactiontime="+12" />
                    <RELAYPOSITION number="3" athleteid="151685" reactiontime="+8" />
                    <RELAYPOSITION number="4" athleteid="213133" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="27" place="13" lane="3" heat="4" swimtime="00:01:34.98" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.82" />
                    <SPLIT distance="50" swimtime="00:00:22.48" />
                    <SPLIT distance="75" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:00:44.84" />
                    <SPLIT distance="125" swimtime="00:00:56.58" />
                    <SPLIT distance="150" swimtime="00:01:09.64" />
                    <SPLIT distance="175" swimtime="00:01:21.85" />
                    <SPLIT distance="200" swimtime="00:01:34.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="151685" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="213133" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="100989" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="129491" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="8" place="11" lane="7" heat="1" swimtime="00:03:40.28" reactiontime="+71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                    <SPLIT distance="75" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:00:54.12" />
                    <SPLIT distance="125" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:20.45" />
                    <SPLIT distance="175" swimtime="00:01:34.85" />
                    <SPLIT distance="200" swimtime="00:01:49.27" />
                    <SPLIT distance="225" swimtime="00:02:01.58" />
                    <SPLIT distance="250" swimtime="00:02:15.66" />
                    <SPLIT distance="275" swimtime="00:02:30.24" />
                    <SPLIT distance="300" swimtime="00:02:45.09" />
                    <SPLIT distance="325" swimtime="00:02:57.35" />
                    <SPLIT distance="350" swimtime="00:03:11.52" />
                    <SPLIT distance="375" swimtime="00:03:26.05" />
                    <SPLIT distance="400" swimtime="00:03:40.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100989" reactiontime="+71" />
                    <RELAYPOSITION number="2" athleteid="101305" reactiontime="+48" />
                    <RELAYPOSITION number="3" athleteid="101068" reactiontime="+45" />
                    <RELAYPOSITION number="4" athleteid="129491" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="47" place="14" lane="1" heat="2" swimtime="00:04:05.26" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="75" swimtime="00:00:46.06" />
                    <SPLIT distance="100" swimtime="00:01:01.82" />
                    <SPLIT distance="125" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:01:33.71" />
                    <SPLIT distance="175" swimtime="00:01:52.10" />
                    <SPLIT distance="200" swimtime="00:02:10.92" />
                    <SPLIT distance="225" swimtime="00:02:23.53" />
                    <SPLIT distance="250" swimtime="00:02:38.92" />
                    <SPLIT distance="275" swimtime="00:02:54.93" />
                    <SPLIT distance="300" swimtime="00:03:11.23" />
                    <SPLIT distance="325" swimtime="00:03:23.19" />
                    <SPLIT distance="350" swimtime="00:03:36.79" />
                    <SPLIT distance="375" swimtime="00:03:51.01" />
                    <SPLIT distance="400" swimtime="00:04:05.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="210408" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="151671" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="214617" reactiontime="+36" />
                    <RELAYPOSITION number="4" athleteid="100989" reactiontime="+54" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="17" place="11" lane="6" heat="2" swimtime="00:08:07.50" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="75" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:00:58.61" />
                    <SPLIT distance="125" swimtime="00:01:14.32" />
                    <SPLIT distance="150" swimtime="00:01:30.84" />
                    <SPLIT distance="175" swimtime="00:01:47.05" />
                    <SPLIT distance="200" swimtime="00:02:03.02" />
                    <SPLIT distance="225" swimtime="00:02:16.04" />
                    <SPLIT distance="250" swimtime="00:02:30.57" />
                    <SPLIT distance="275" swimtime="00:02:45.60" />
                    <SPLIT distance="300" swimtime="00:03:01.00" />
                    <SPLIT distance="325" swimtime="00:03:16.51" />
                    <SPLIT distance="350" swimtime="00:03:32.53" />
                    <SPLIT distance="375" swimtime="00:03:48.55" />
                    <SPLIT distance="400" swimtime="00:04:03.90" />
                    <SPLIT distance="425" swimtime="00:04:16.01" />
                    <SPLIT distance="450" swimtime="00:04:30.20" />
                    <SPLIT distance="475" swimtime="00:04:44.69" />
                    <SPLIT distance="500" swimtime="00:04:59.80" />
                    <SPLIT distance="525" swimtime="00:05:15.20" />
                    <SPLIT distance="550" swimtime="00:05:30.90" />
                    <SPLIT distance="575" swimtime="00:05:47.23" />
                    <SPLIT distance="600" swimtime="00:06:02.93" />
                    <SPLIT distance="625" swimtime="00:06:15.96" />
                    <SPLIT distance="650" swimtime="00:06:31.08" />
                    <SPLIT distance="675" swimtime="00:06:46.68" />
                    <SPLIT distance="700" swimtime="00:07:02.67" />
                    <SPLIT distance="725" swimtime="00:07:18.82" />
                    <SPLIT distance="750" swimtime="00:07:35.20" />
                    <SPLIT distance="775" swimtime="00:07:51.61" />
                    <SPLIT distance="800" swimtime="00:08:07.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="210412" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="129491" reactiontime="+43" />
                    <RELAYPOSITION number="3" athleteid="100989" reactiontime="+46" />
                    <RELAYPOSITION number="4" athleteid="151671" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="25" place="9" lane="3" heat="2" swimtime="00:01:40.36" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.10" />
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                    <SPLIT distance="75" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:00:49.61" />
                    <SPLIT distance="125" swimtime="00:01:02.08" />
                    <SPLIT distance="150" swimtime="00:01:15.26" />
                    <SPLIT distance="175" swimtime="00:01:27.29" />
                    <SPLIT distance="200" swimtime="00:01:40.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100989" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="101305" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="129491" reactiontime="+30" />
                    <RELAYPOSITION number="4" athleteid="101068" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="34" place="12" lane="6" heat="1" swimtime="00:01:52.61" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                    <SPLIT distance="75" swimtime="00:00:41.87" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                    <SPLIT distance="125" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:26.39" />
                    <SPLIT distance="175" swimtime="00:01:38.91" />
                    <SPLIT distance="200" swimtime="00:01:52.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101305" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="151671" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="101068" reactiontime="+42" />
                    <RELAYPOSITION number="4" athleteid="214616" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="11" place="14" lane="3" heat="2" swimtime="00:01:42.05" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:00:55.41" />
                    <SPLIT distance="125" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:21.34" />
                    <SPLIT distance="175" swimtime="00:01:31.13" />
                    <SPLIT distance="200" swimtime="00:01:42.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101305" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="105413" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="100989" reactiontime="+38" />
                    <RELAYPOSITION number="4" athleteid="165123" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Hong Kong, China">
              <RESULTS>
                <RESULT eventid="35" place="11" lane="4" heat="1" swimtime="00:01:34.74" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:00:51.81" />
                    <SPLIT distance="125" swimtime="00:01:01.93" />
                    <SPLIT distance="150" swimtime="00:01:14.40" />
                    <SPLIT distance="175" swimtime="00:01:23.98" />
                    <SPLIT distance="200" swimtime="00:01:34.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213133" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="105413" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="151685" reactiontime="+14" />
                    <RELAYPOSITION number="4" athleteid="165123" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Honduras" shortname="HON" code="HON" nation="HON" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="145120" lastname="HORREGO" firstname="Julio" gender="M" birthdate="1998-10-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.80" eventid="16" heat="4" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.38" eventid="41" heat="5" lane="3">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="34" lane="4" heat="4" heatid="40016" swimtime="00:00:59.22" reactiontime="+68" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="75" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:00:59.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="39" lane="3" heat="5" heatid="50041" swimtime="00:00:27.71" reactiontime="+63" points="729">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130156" lastname="VASQUEZ" firstname="Carlos" gender="M" birthdate="2000-06-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.91" eventid="39" heat="3" lane="3">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:01:58.41" eventid="21" heat="4" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="38" lane="3" heat="3" heatid="30039" swimtime="00:00:53.36" reactiontime="+61" points="717">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                    <SPLIT distance="75" swimtime="00:00:39.15" />
                    <SPLIT distance="100" swimtime="00:00:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="22" lane="8" heat="4" heatid="40021" swimtime="00:01:58.63" reactiontime="+64" points="759">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.05" />
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="75" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:00:55.75" />
                    <SPLIT distance="125" swimtime="00:01:10.84" />
                    <SPLIT distance="150" swimtime="00:01:26.24" />
                    <SPLIT distance="175" swimtime="00:01:42.14" />
                    <SPLIT distance="200" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100488" lastname="AVILA MANCIA" firstname="Julimar" gender="F" birthdate="1997-01-21">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.18" eventid="38" heat="1" lane="7">
                  <MEETINFO date="2022-04-22" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.68" eventid="43" heat="2" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="26" lane="7" heat="1" heatid="10038" swimtime="00:01:01.43" reactiontime="+68" points="701">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="75" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="28" lane="7" heat="2" heatid="20043" swimtime="00:02:04.28" reactiontime="+71" points="699">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                    <SPLIT distance="75" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:01:00.26" />
                    <SPLIT distance="125" swimtime="00:01:16.12" />
                    <SPLIT distance="150" swimtime="00:01:32.25" />
                    <SPLIT distance="175" swimtime="00:01:48.49" />
                    <SPLIT distance="200" swimtime="00:02:04.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Hungary" shortname="HUN" code="HUN" nation="HUN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="166325" lastname="SZABO" firstname="Szebasztian" gender="M" birthdate="1996-03-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.68" eventid="39" heat="6" lane="3">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:47.14" eventid="14" heat="10" lane="8">
                  <MEETINFO date="2021-10-08" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.75" eventid="5" heat="10" lane="4">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:20.72" eventid="31" heat="11" lane="5">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="-1" lane="3" heat="6" heatid="60039" swimtime="NT" status="DNS" />
                <RESULT eventid="14" place="18" lane="8" heat="10" heatid="100014" swimtime="00:00:47.09" reactiontime="+61" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.53" />
                    <SPLIT distance="50" swimtime="00:00:22.56" />
                    <SPLIT distance="75" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:00:47.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="105" place="3" lane="4" heat="1" heatid="10105" swimtime="00:00:21.98" reactiontime="+58" points="968">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.91" />
                    <SPLIT distance="50" swimtime="00:00:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="3" lane="4" heat="10" heatid="100005" swimtime="00:00:22.07" reactiontime="+58" points="957">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.02" />
                    <SPLIT distance="50" swimtime="00:00:22.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="1" lane="5" heat="2" heatid="20205" swimtime="00:00:21.90" reactiontime="+57" points="979">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.87" />
                    <SPLIT distance="50" swimtime="00:00:21.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="131" place="4" lane="3" heat="1" heatid="10131" swimtime="00:00:20.84" reactiontime="+59" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.91" />
                    <SPLIT distance="50" swimtime="00:00:20.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="6" lane="5" heat="11" heatid="110031" swimtime="00:00:21.00" reactiontime="+64" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.08" />
                    <SPLIT distance="50" swimtime="00:00:21.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="3" lane="6" heat="2" heatid="20231" swimtime="00:00:20.83" reactiontime="+57" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.87" />
                    <SPLIT distance="50" swimtime="00:00:20.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101670" lastname="JAKABOS" firstname="Zsuzsanna" gender="F" birthdate="1989-04-03">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.67" eventid="20" heat="3" lane="6">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.36" eventid="43" heat="3" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.94" eventid="6" heat="5" lane="3">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:04:30.38" eventid="36" heat="3" lane="3">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="13" lane="6" heat="3" heatid="30020" swimtime="00:02:07.08" reactiontime="+74" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="75" swimtime="00:00:44.86" />
                    <SPLIT distance="100" swimtime="00:01:01.01" />
                    <SPLIT distance="125" swimtime="00:01:17.32" />
                    <SPLIT distance="150" swimtime="00:01:33.76" />
                    <SPLIT distance="175" swimtime="00:01:50.33" />
                    <SPLIT distance="200" swimtime="00:02:07.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="-1" lane="2" heat="3" heatid="30043" swimtime="NT" status="DNS" />
                <RESULT eventid="6" place="16" lane="3" heat="5" heatid="50006" swimtime="00:02:09.63" reactiontime="+75" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:44.79" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="125" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:01:38.78" />
                    <SPLIT distance="175" swimtime="00:01:55.16" />
                    <SPLIT distance="200" swimtime="00:02:09.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="5" lane="6" heat="1" heatid="10136" swimtime="00:04:32.10" reactiontime="+74" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="75" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="125" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:01:37.70" />
                    <SPLIT distance="175" swimtime="00:01:54.94" />
                    <SPLIT distance="200" swimtime="00:02:11.83" />
                    <SPLIT distance="225" swimtime="00:02:31.48" />
                    <SPLIT distance="250" swimtime="00:02:51.37" />
                    <SPLIT distance="275" swimtime="00:03:11.09" />
                    <SPLIT distance="300" swimtime="00:03:31.23" />
                    <SPLIT distance="325" swimtime="00:03:47.05" />
                    <SPLIT distance="350" swimtime="00:04:02.05" />
                    <SPLIT distance="375" swimtime="00:04:17.31" />
                    <SPLIT distance="400" swimtime="00:04:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="4" lane="3" heat="3" heatid="30036" swimtime="00:04:31.36" reactiontime="+74" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="75" swimtime="00:00:45.87" />
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                    <SPLIT distance="125" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:01:36.62" />
                    <SPLIT distance="175" swimtime="00:01:53.56" />
                    <SPLIT distance="200" swimtime="00:02:10.17" />
                    <SPLIT distance="225" swimtime="00:02:29.65" />
                    <SPLIT distance="250" swimtime="00:02:49.46" />
                    <SPLIT distance="275" swimtime="00:03:09.43" />
                    <SPLIT distance="300" swimtime="00:03:29.18" />
                    <SPLIT distance="325" swimtime="00:03:45.49" />
                    <SPLIT distance="350" swimtime="00:04:01.03" />
                    <SPLIT distance="375" swimtime="00:04:16.48" />
                    <SPLIT distance="400" swimtime="00:04:31.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="India" shortname="IND" code="IND" nation="IND" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="213832" lastname="SRIDHAR" firstname="Siva" gender="M" birthdate="2000-11-07">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="7" heat="1" lane="7" />
                <ENTRY entrytime="NT" eventid="23" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="30" lane="7" heat="1" heatid="10007" swimtime="00:01:59.80" reactiontime="+68" points="766">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.51" />
                    <SPLIT distance="50" swimtime="00:00:25.28" />
                    <SPLIT distance="75" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:00:54.57" />
                    <SPLIT distance="125" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:29.80" />
                    <SPLIT distance="175" swimtime="00:01:45.30" />
                    <SPLIT distance="200" swimtime="00:01:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="33" lane="5" heat="1" heatid="10023" swimtime="00:00:56.80" reactiontime="+67" points="653">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.47" />
                    <SPLIT distance="50" swimtime="00:00:25.40" />
                    <SPLIT distance="75" swimtime="00:00:42.37" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213831" lastname="ARORA" firstname="Chahat" gender="F" birthdate="1997-07-17">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="15" heat="1" lane="6" />
                <ENTRY entrytime="NT" eventid="40" heat="2" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="42" lane="6" heat="1" heatid="10015" swimtime="00:01:13.13" reactiontime="+67" points="620">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.94" />
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="75" swimtime="00:00:53.19" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="31" lane="1" heat="2" heatid="20040" swimtime="00:00:32.91" reactiontime="+57" points="653">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.16" />
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Islamic Rep. of Iran" shortname="IRI" code="IRI" nation="IRI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="179236" lastname="AFGHARI" firstname="Mehrshad" gender="M" birthdate="2001-11-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.87" eventid="39" heat="4" lane="5">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="36" lane="5" heat="4" heatid="40039" swimtime="00:00:52.95" reactiontime="+68" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:24.81" />
                    <SPLIT distance="75" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:00:52.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140761" lastname="GHOLAMPOUR" firstname="Sina" gender="M" birthdate="1999-09-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.60" eventid="14" heat="6" lane="5">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.26" eventid="31" heat="6" lane="6">
                  <MEETINFO date="2021-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="-1" lane="5" heat="6" heatid="60014" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="-1" lane="6" heat="6" heatid="60031" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Iraq" shortname="IRQ" code="IRQ" nation="IRQ" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198120" lastname="AL-HASANI" firstname="Ahmed Alaa  Jabbar" gender="M" birthdate="2006-03-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:07.98" eventid="16" heat="1" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.81" eventid="14" heat="3" lane="2">
                  <MEETINFO date="2021-10-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="56" lane="4" heat="1" heatid="10016" swimtime="00:01:06.77" reactiontime="+67" points="567">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                    <SPLIT distance="75" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:06.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="63" lane="2" heat="3" heatid="30014" swimtime="00:00:51.96" reactiontime="+67" points="642">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:24.97" />
                    <SPLIT distance="75" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:00:51.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Iceland" shortname="ISL" code="ISL" nation="ISL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="100751" lastname="MCKEE" firstname="Anton " gender="M" birthdate="1993-12-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.53" eventid="16" heat="6" lane="7">
                  <MEETINFO date="2021-11-14" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.54" eventid="29" heat="5" lane="3">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.91" eventid="41" heat="6" lane="3">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="18" lane="7" heat="6" heatid="60016" swimtime="00:00:58.01" reactiontime="+62" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="75" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:00:58.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="10" lane="3" heat="5" heatid="50029" swimtime="00:02:04.99" reactiontime="+63" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.85" />
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="75" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:00:59.88" />
                    <SPLIT distance="125" swimtime="00:01:15.83" />
                    <SPLIT distance="150" swimtime="00:01:31.99" />
                    <SPLIT distance="175" swimtime="00:01:48.42" />
                    <SPLIT distance="200" swimtime="00:02:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="-1" lane="3" heat="6" heatid="60041" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164729" lastname="JÓRUNNARDÓTTIR" firstname="Snæfríður Sól" gender="F" birthdate="2000-10-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.99" eventid="13" heat="6" lane="6">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.47" eventid="43" heat="3" lane="7">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="15" lane="6" heat="6" heatid="60013" swimtime="00:00:53.21" reactiontime="+68" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.37" />
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                    <SPLIT distance="75" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="15" lane="8" heat="2" heatid="20213" swimtime="00:00:53.19" reactiontime="+69" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.72" />
                    <SPLIT distance="75" swimtime="00:00:39.41" />
                    <SPLIT distance="100" swimtime="00:00:53.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="11" lane="7" heat="3" heatid="30043" swimtime="00:01:55.34" reactiontime="+71" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="75" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:00:57.14" />
                    <SPLIT distance="125" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:26.53" />
                    <SPLIT distance="175" swimtime="00:01:41.14" />
                    <SPLIT distance="200" swimtime="00:01:55.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Israel" shortname="ISR" code="ISR" nation="ISR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="144949" lastname="CHERUTI" firstname="Meiron Amir" gender="M" birthdate="1997-10-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.49" eventid="14" heat="6" lane="4">
                  <MEETINFO date="2021-09-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.44" eventid="19" heat="2" lane="6">
                  <MEETINFO date="2022-05-12" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.58" eventid="5" heat="5" lane="7">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.95" eventid="31" heat="7" lane="6">
                  <MEETINFO date="2022-05-11" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="42" lane="4" heat="6" heatid="60014" swimtime="00:00:48.20" reactiontime="+65" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.57" />
                    <SPLIT distance="50" swimtime="00:00:22.38" />
                    <SPLIT distance="75" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:00:48.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="-1" lane="6" heat="2" heatid="20019" swimtime="00:00:24.12" status="DSQ" reactiontime="+62" />
                <RESULT eventid="5" place="26" lane="7" heat="5" heatid="50005" swimtime="00:00:22.90" reactiontime="+65" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.31" />
                    <SPLIT distance="50" swimtime="00:00:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="18" lane="6" heat="7" heatid="70031" swimtime="00:00:21.33" reactiontime="+63" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.15" />
                    <SPLIT distance="50" swimtime="00:00:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="331" place="20" lane="4" heat="1" heatid="10331" swimtime="00:00:21.45" reactiontime="+63" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100840" lastname="TOUMARKIN" firstname="Yakov" gender="M" birthdate="1992-02-15">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.55" eventid="46" heat="4" lane="7">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.97" eventid="7" heat="4" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.17" eventid="23" heat="5" lane="2">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="13" lane="7" heat="4" heatid="40046" swimtime="00:01:53.03" reactiontime="+60" points="816">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                    <SPLIT distance="75" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:00:55.32" />
                    <SPLIT distance="125" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:24.47" />
                    <SPLIT distance="175" swimtime="00:01:39.00" />
                    <SPLIT distance="200" swimtime="00:01:53.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="16" lane="2" heat="4" heatid="40007" swimtime="00:01:54.95" reactiontime="+65" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="75" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:00:53.85" />
                    <SPLIT distance="125" swimtime="00:01:10.13" />
                    <SPLIT distance="150" swimtime="00:01:26.87" />
                    <SPLIT distance="175" swimtime="00:01:41.53" />
                    <SPLIT distance="200" swimtime="00:01:54.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="10" lane="2" heat="5" heatid="50023" swimtime="00:00:52.38" reactiontime="+67" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.82" />
                    <SPLIT distance="50" swimtime="00:00:23.75" />
                    <SPLIT distance="75" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:00:52.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="14" lane="2" heat="1" heatid="10223" swimtime="00:00:52.74" reactiontime="+63" points="815">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.64" />
                    <SPLIT distance="75" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:00:52.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Virgin Islands, US" shortname="ISV" code="ISV" nation="ISV" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="182690" lastname="WILSON" firstname="Maximillian" gender="M" birthdate="2004-04-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.21" eventid="3" heat="3" lane="8">
                  <MEETINFO date="2021-10-31" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.18" eventid="19" heat="2" lane="4">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="32" lane="8" heat="3" heatid="30003" swimtime="00:00:53.23" reactiontime="+58" points="748">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:25.38" />
                    <SPLIT distance="75" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:00:53.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="30" lane="4" heat="2" heatid="20019" swimtime="00:00:24.31" reactiontime="+57" points="763">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:24.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121632" lastname="SANES" firstname="Adriel " gender="M" birthdate="1998-10-27">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.71" eventid="29" heat="2" lane="7">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.25" eventid="41" heat="4" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="29" place="27" lane="7" heat="2" heatid="20029" swimtime="00:02:12.69" reactiontime="+65" points="742">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.23" />
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="75" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="125" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:01:37.45" />
                    <SPLIT distance="175" swimtime="00:01:54.90" />
                    <SPLIT distance="200" swimtime="00:02:12.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="40" lane="2" heat="4" heatid="40041" swimtime="00:00:27.76" reactiontime="+64" points="726">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.50" />
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150470" lastname="KUIPERS" firstname="Natalia Jean" gender="F" birthdate="2002-06-13">
              <ENTRIES>
                <ENTRY entrytime="00:04:26.48" eventid="1" heat="1" lane="3">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:09:32.24" eventid="12" heat="1" lane="7">
                  <MEETINFO date="2022-07-09" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="26" lane="3" heat="1" heatid="10001" swimtime="00:04:26.11" reactiontime="+73" points="679">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="75" swimtime="00:00:45.62" />
                    <SPLIT distance="100" swimtime="00:01:01.80" />
                    <SPLIT distance="125" swimtime="00:01:18.23" />
                    <SPLIT distance="150" swimtime="00:01:34.97" />
                    <SPLIT distance="175" swimtime="00:01:51.62" />
                    <SPLIT distance="200" swimtime="00:02:08.72" />
                    <SPLIT distance="225" swimtime="00:02:25.79" />
                    <SPLIT distance="250" swimtime="00:02:43.02" />
                    <SPLIT distance="275" swimtime="00:03:00.25" />
                    <SPLIT distance="300" swimtime="00:03:17.50" />
                    <SPLIT distance="325" swimtime="00:03:34.74" />
                    <SPLIT distance="350" swimtime="00:03:52.27" />
                    <SPLIT distance="375" swimtime="00:04:09.54" />
                    <SPLIT distance="400" swimtime="00:04:26.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="20" lane="7" heat="1" heatid="10012" swimtime="00:09:03.17" reactiontime="+74" points="687">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="75" swimtime="00:00:46.68" />
                    <SPLIT distance="100" swimtime="00:01:03.52" />
                    <SPLIT distance="125" swimtime="00:01:20.27" />
                    <SPLIT distance="150" swimtime="00:01:37.16" />
                    <SPLIT distance="175" swimtime="00:01:53.91" />
                    <SPLIT distance="200" swimtime="00:02:10.80" />
                    <SPLIT distance="225" swimtime="00:02:27.64" />
                    <SPLIT distance="250" swimtime="00:02:44.64" />
                    <SPLIT distance="275" swimtime="00:03:01.59" />
                    <SPLIT distance="300" swimtime="00:03:18.83" />
                    <SPLIT distance="325" swimtime="00:03:35.91" />
                    <SPLIT distance="350" swimtime="00:03:53.19" />
                    <SPLIT distance="375" swimtime="00:04:10.41" />
                    <SPLIT distance="400" swimtime="00:04:27.76" />
                    <SPLIT distance="425" swimtime="00:04:44.88" />
                    <SPLIT distance="450" swimtime="00:05:02.13" />
                    <SPLIT distance="475" swimtime="00:05:19.33" />
                    <SPLIT distance="500" swimtime="00:05:36.60" />
                    <SPLIT distance="525" swimtime="00:05:53.83" />
                    <SPLIT distance="550" swimtime="00:06:11.06" />
                    <SPLIT distance="575" swimtime="00:06:28.39" />
                    <SPLIT distance="600" swimtime="00:06:45.62" />
                    <SPLIT distance="625" swimtime="00:07:02.98" />
                    <SPLIT distance="650" swimtime="00:07:20.25" />
                    <SPLIT distance="675" swimtime="00:07:37.49" />
                    <SPLIT distance="700" swimtime="00:07:54.76" />
                    <SPLIT distance="725" swimtime="00:08:12.12" />
                    <SPLIT distance="750" swimtime="00:08:29.37" />
                    <SPLIT distance="775" swimtime="00:08:46.65" />
                    <SPLIT distance="800" swimtime="00:09:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Italy" shortname="ITA" code="ITA" nation="ITA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154842" lastname="MORA" firstname="Lorenzo" gender="M" birthdate="1998-09-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.37" eventid="3" heat="5" lane="4">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:01:48.72" eventid="46" heat="4" lane="5">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.90" eventid="19" heat="5" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="2" lane="3" heat="1" heatid="10103" swimtime="00:00:49.04" reactiontime="+52" points="957">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:24.04" />
                    <SPLIT distance="75" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="7" lane="4" heat="5" heatid="50003" swimtime="00:00:50.18" reactiontime="+61" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:24.22" />
                    <SPLIT distance="75" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:00:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="3" lane="6" heat="2" heatid="20203" swimtime="00:00:49.57" reactiontime="+55" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.69" />
                    <SPLIT distance="50" swimtime="00:00:24.16" />
                    <SPLIT distance="75" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:00:49.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="146" place="3" lane="6" heat="1" heatid="10146" swimtime="00:01:48.45" reactiontime="+56" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                    <SPLIT distance="75" swimtime="00:00:40.11" />
                    <SPLIT distance="100" swimtime="00:00:54.13" />
                    <SPLIT distance="125" swimtime="00:01:07.76" />
                    <SPLIT distance="150" swimtime="00:01:21.70" />
                    <SPLIT distance="175" swimtime="00:01:35.02" />
                    <SPLIT distance="200" swimtime="00:01:48.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="4" lane="5" heat="4" heatid="40046" swimtime="00:01:49.79" reactiontime="+60" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                    <SPLIT distance="50" swimtime="00:00:26.12" />
                    <SPLIT distance="75" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:00:54.12" />
                    <SPLIT distance="125" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:21.96" />
                    <SPLIT distance="175" swimtime="00:01:35.89" />
                    <SPLIT distance="200" swimtime="00:01:49.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="4" lane="7" heat="1" heatid="10119" swimtime="00:00:22.81" reactiontime="+53" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.06" />
                    <SPLIT distance="50" swimtime="00:00:22.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="5" lane="5" heat="5" heatid="50019" swimtime="00:00:23.09" reactiontime="+55" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:23.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="5" lane="3" heat="2" heatid="20219" swimtime="00:00:22.90" reactiontime="+55" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.20" />
                    <SPLIT distance="50" swimtime="00:00:22.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124772" lastname="MARTINENGHI" firstname="Nicolò" gender="M" birthdate="1999-08-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.63" eventid="16" heat="7" lane="4">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:25.37" eventid="41" heat="9" lane="4">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="2" lane="4" heat="1" heatid="10116" swimtime="00:00:56.07" reactiontime="+62" points="958">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:26.36" />
                    <SPLIT distance="75" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:00:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="1" lane="4" heat="7" heatid="70016" swimtime="00:00:56.60" reactiontime="+63" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                    <SPLIT distance="75" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:00:56.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="1" lane="4" heat="2" heatid="20216" swimtime="00:00:56.01" reactiontime="+62" points="961">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                    <SPLIT distance="75" swimtime="00:00:40.96" />
                    <SPLIT distance="100" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="2" lane="4" heat="1" heatid="10141" swimtime="00:00:25.42" reactiontime="+61" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:25.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="1" lane="4" heat="9" heatid="90041" swimtime="00:00:25.71" reactiontime="+63" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:25.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="1" lane="4" heat="2" heatid="20241" swimtime="00:00:25.60" reactiontime="+62" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198800" lastname="CERASUOLO" firstname="Simone" gender="M" birthdate="2003-06-22">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.80" eventid="16" heat="8" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:25.78" eventid="41" heat="9" lane="5">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="6" lane="2" heat="1" heatid="10116" swimtime="00:00:56.99" reactiontime="+63" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                    <SPLIT distance="75" swimtime="00:00:41.74" />
                    <SPLIT distance="100" swimtime="00:00:56.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="9" lane="3" heat="8" heatid="80016" swimtime="00:00:57.24" reactiontime="+64" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.95" />
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                    <SPLIT distance="75" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:00:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="5" lane="2" heat="2" heatid="20216" swimtime="00:00:56.71" reactiontime="+63" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.79" />
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                    <SPLIT distance="75" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:00:56.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="3" lane="3" heat="1" heatid="10141" swimtime="00:00:25.68" reactiontime="+65" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:25.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="7" lane="5" heat="9" heatid="90041" swimtime="00:00:26.16" reactiontime="+65" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="3" lane="6" heat="2" heatid="20241" swimtime="00:00:25.66" reactiontime="+62" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:25.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102367" lastname="RIVOLTA" firstname="Matteo" gender="M" birthdate="1991-11-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.64" eventid="39" heat="7" lane="4">
                  <MEETINFO date="2021-11-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.02" eventid="5" heat="10" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="5" lane="5" heat="1" heatid="10139" swimtime="00:00:49.32" reactiontime="+68" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.43" />
                    <SPLIT distance="50" swimtime="00:00:22.72" />
                    <SPLIT distance="75" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:00:49.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="2" lane="4" heat="7" heatid="70039" swimtime="00:00:49.43" reactiontime="+65" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:22.76" />
                    <SPLIT distance="75" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:00:49.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="2" lane="4" heat="1" heatid="10239" swimtime="00:00:49.07" reactiontime="+66" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.38" />
                    <SPLIT distance="50" swimtime="00:00:22.81" />
                    <SPLIT distance="75" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="8" lane="5" heat="10" heatid="100005" swimtime="00:00:22.32" reactiontime="+67" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.30" />
                    <SPLIT distance="50" swimtime="00:00:22.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="-1" lane="2" heat="2" heatid="20205" swimtime="00:00:22.56" status="DSQ" reactiontime="+65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124771" lastname="MIRESSI" firstname="Alessandro" gender="M" birthdate="1998-10-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:45.57" eventid="14" heat="10" lane="4">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.20" eventid="31" heat="10" lane="2">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="3" lane="6" heat="1" heatid="10114" swimtime="00:00:45.57" reactiontime="+68" points="952">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.73" />
                    <SPLIT distance="75" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="5" lane="4" heat="10" heatid="100014" swimtime="00:00:46.22" reactiontime="+68" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.41" />
                    <SPLIT distance="50" swimtime="00:00:22.04" />
                    <SPLIT distance="75" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:00:46.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="4" lane="3" heat="2" heatid="20214" swimtime="00:00:45.74" reactiontime="+69" points="942">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.29" />
                    <SPLIT distance="50" swimtime="00:00:21.90" />
                    <SPLIT distance="75" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:00:45.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="12" lane="2" heat="10" heatid="100031" swimtime="00:00:21.17" reactiontime="+67" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.22" />
                    <SPLIT distance="50" swimtime="00:00:21.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="13" lane="7" heat="2" heatid="20231" swimtime="00:00:21.13" reactiontime="+68" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.11" />
                    <SPLIT distance="50" swimtime="00:00:21.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149646" lastname="CECCON" firstname="Thomas" gender="M" birthdate="2001-01-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.15" eventid="14" heat="11" lane="5">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.19" eventid="5" heat="9" lane="5">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.40" eventid="23" heat="5" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="5" lane="7" heat="1" heatid="10114" swimtime="00:00:45.72" reactiontime="+68" points="943">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.29" />
                    <SPLIT distance="50" swimtime="00:00:21.97" />
                    <SPLIT distance="75" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="7" lane="5" heat="11" heatid="110014" swimtime="00:00:46.41" reactiontime="+68" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:22.09" />
                    <SPLIT distance="75" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="6" lane="6" heat="2" heatid="20214" swimtime="00:00:46.13" reactiontime="+68" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.34" />
                    <SPLIT distance="50" swimtime="00:00:21.92" />
                    <SPLIT distance="75" swimtime="00:00:34.03" />
                    <SPLIT distance="100" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="19" lane="5" heat="9" heatid="90005" swimtime="00:00:22.57" reactiontime="+68" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.20" />
                    <SPLIT distance="50" swimtime="00:00:22.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="1" lane="2" heat="1" heatid="10123" swimtime="00:00:50.97" reactiontime="+67" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.37" />
                    <SPLIT distance="50" swimtime="00:00:22.77" />
                    <SPLIT distance="75" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:00:50.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="6" lane="5" heat="5" heatid="50023" swimtime="00:00:52.12" reactiontime="+69" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.54" />
                    <SPLIT distance="50" swimtime="00:00:23.34" />
                    <SPLIT distance="75" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:00:52.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="5" lane="3" heat="1" heatid="10223" swimtime="00:00:51.60" reactiontime="+67" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.36" />
                    <SPLIT distance="50" swimtime="00:00:23.21" />
                    <SPLIT distance="75" swimtime="00:00:38.57" />
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101853" lastname="PALTRINIERI" firstname="Gregorio" gender="M" birthdate="1994-09-05">
              <ENTRIES>
                <ENTRY entrytime="00:14:13.07" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:07:27.94" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="1" lane="4" heat="5" heatid="30110" swimtime="00:14:16.88" reactiontime="+78" points="965">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                    <SPLIT distance="75" swimtime="00:00:40.16" />
                    <SPLIT distance="100" swimtime="00:00:54.10" />
                    <SPLIT distance="125" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:22.35" />
                    <SPLIT distance="175" swimtime="00:01:36.54" />
                    <SPLIT distance="200" swimtime="00:01:50.90" />
                    <SPLIT distance="225" swimtime="00:02:05.27" />
                    <SPLIT distance="250" swimtime="00:02:19.69" />
                    <SPLIT distance="275" swimtime="00:02:33.99" />
                    <SPLIT distance="300" swimtime="00:02:48.41" />
                    <SPLIT distance="325" swimtime="00:03:02.71" />
                    <SPLIT distance="350" swimtime="00:03:17.04" />
                    <SPLIT distance="375" swimtime="00:03:31.32" />
                    <SPLIT distance="400" swimtime="00:03:45.69" />
                    <SPLIT distance="425" swimtime="00:04:00.14" />
                    <SPLIT distance="450" swimtime="00:04:14.71" />
                    <SPLIT distance="475" swimtime="00:04:29.07" />
                    <SPLIT distance="500" swimtime="00:04:43.61" />
                    <SPLIT distance="525" swimtime="00:04:57.95" />
                    <SPLIT distance="550" swimtime="00:05:12.44" />
                    <SPLIT distance="575" swimtime="00:05:26.72" />
                    <SPLIT distance="600" swimtime="00:05:41.13" />
                    <SPLIT distance="625" swimtime="00:05:55.44" />
                    <SPLIT distance="650" swimtime="00:06:09.76" />
                    <SPLIT distance="675" swimtime="00:06:24.15" />
                    <SPLIT distance="700" swimtime="00:06:38.54" />
                    <SPLIT distance="725" swimtime="00:06:52.97" />
                    <SPLIT distance="750" swimtime="00:07:07.31" />
                    <SPLIT distance="775" swimtime="00:07:21.72" />
                    <SPLIT distance="800" swimtime="00:07:35.98" />
                    <SPLIT distance="825" swimtime="00:07:50.43" />
                    <SPLIT distance="850" swimtime="00:08:04.76" />
                    <SPLIT distance="875" swimtime="00:08:19.12" />
                    <SPLIT distance="900" swimtime="00:08:33.54" />
                    <SPLIT distance="925" swimtime="00:08:47.87" />
                    <SPLIT distance="950" swimtime="00:09:02.23" />
                    <SPLIT distance="975" swimtime="00:09:16.59" />
                    <SPLIT distance="1000" swimtime="00:09:30.83" />
                    <SPLIT distance="1025" swimtime="00:09:45.18" />
                    <SPLIT distance="1050" swimtime="00:09:59.43" />
                    <SPLIT distance="1075" swimtime="00:10:13.91" />
                    <SPLIT distance="1100" swimtime="00:10:28.20" />
                    <SPLIT distance="1125" swimtime="00:10:42.69" />
                    <SPLIT distance="1150" swimtime="00:10:57.01" />
                    <SPLIT distance="1175" swimtime="00:11:11.38" />
                    <SPLIT distance="1200" swimtime="00:11:25.65" />
                    <SPLIT distance="1225" swimtime="00:11:39.65" />
                    <SPLIT distance="1250" swimtime="00:11:53.87" />
                    <SPLIT distance="1275" swimtime="00:12:08.15" />
                    <SPLIT distance="1300" swimtime="00:12:22.33" />
                    <SPLIT distance="1325" swimtime="00:12:36.53" />
                    <SPLIT distance="1350" swimtime="00:12:50.77" />
                    <SPLIT distance="1375" swimtime="00:13:05.20" />
                    <SPLIT distance="1400" swimtime="00:13:19.64" />
                    <SPLIT distance="1425" swimtime="00:13:34.26" />
                    <SPLIT distance="1450" swimtime="00:13:48.80" />
                    <SPLIT distance="1475" swimtime="00:14:03.21" />
                    <SPLIT distance="1500" swimtime="00:14:16.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="1" lane="4" heat="5" heatid="30142" swimtime="00:07:29.99" reactiontime="+78" points="956">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                    <SPLIT distance="75" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:00:53.98" />
                    <SPLIT distance="125" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:22.48" />
                    <SPLIT distance="175" swimtime="00:01:36.77" />
                    <SPLIT distance="200" swimtime="00:01:51.15" />
                    <SPLIT distance="225" swimtime="00:02:05.55" />
                    <SPLIT distance="250" swimtime="00:02:19.87" />
                    <SPLIT distance="275" swimtime="00:02:34.20" />
                    <SPLIT distance="300" swimtime="00:02:48.60" />
                    <SPLIT distance="325" swimtime="00:03:02.94" />
                    <SPLIT distance="350" swimtime="00:03:17.28" />
                    <SPLIT distance="375" swimtime="00:03:31.50" />
                    <SPLIT distance="400" swimtime="00:03:45.81" />
                    <SPLIT distance="425" swimtime="00:03:59.86" />
                    <SPLIT distance="450" swimtime="00:04:13.73" />
                    <SPLIT distance="475" swimtime="00:04:27.66" />
                    <SPLIT distance="500" swimtime="00:04:41.60" />
                    <SPLIT distance="525" swimtime="00:04:55.73" />
                    <SPLIT distance="550" swimtime="00:05:09.82" />
                    <SPLIT distance="575" swimtime="00:05:23.94" />
                    <SPLIT distance="600" swimtime="00:05:38.01" />
                    <SPLIT distance="625" swimtime="00:05:52.08" />
                    <SPLIT distance="650" swimtime="00:06:06.10" />
                    <SPLIT distance="675" swimtime="00:06:20.09" />
                    <SPLIT distance="700" swimtime="00:06:34.14" />
                    <SPLIT distance="725" swimtime="00:06:48.24" />
                    <SPLIT distance="750" swimtime="00:07:02.26" />
                    <SPLIT distance="775" swimtime="00:07:16.35" />
                    <SPLIT distance="800" swimtime="00:07:29.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149648" lastname="RAZZETTI" firstname="Alberto" gender="M" birthdate="1999-06-02">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.06" eventid="21" heat="4" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.54" eventid="7" heat="3" lane="5" />
                <ENTRY entrytime="00:03:59.57" eventid="37" heat="2" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="121" place="4" lane="8" heat="1" heatid="10121" swimtime="00:01:50.12" reactiontime="+70" points="949">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.04" />
                    <SPLIT distance="50" swimtime="00:00:24.67" />
                    <SPLIT distance="75" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:00:52.48" />
                    <SPLIT distance="125" swimtime="00:01:06.58" />
                    <SPLIT distance="150" swimtime="00:01:20.94" />
                    <SPLIT distance="175" swimtime="00:01:35.22" />
                    <SPLIT distance="200" swimtime="00:01:50.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="8" lane="4" heat="4" heatid="40021" swimtime="00:01:50.89" reactiontime="+65" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.36" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:00:53.28" />
                    <SPLIT distance="125" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:21.91" />
                    <SPLIT distance="175" swimtime="00:01:36.29" />
                    <SPLIT distance="200" swimtime="00:01:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="107" place="6" lane="1" heat="1" heatid="10107" swimtime="00:01:51.73" reactiontime="+64" points="944">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.93" />
                    <SPLIT distance="50" swimtime="00:00:23.97" />
                    <SPLIT distance="75" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:00:52.35" />
                    <SPLIT distance="125" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:24.60" />
                    <SPLIT distance="175" swimtime="00:01:38.75" />
                    <SPLIT distance="200" swimtime="00:01:51.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="7" lane="5" heat="3" heatid="30007" swimtime="00:01:52.98" reactiontime="+63" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.90" />
                    <SPLIT distance="50" swimtime="00:00:24.41" />
                    <SPLIT distance="75" swimtime="00:00:39.28" />
                    <SPLIT distance="100" swimtime="00:00:53.18" />
                    <SPLIT distance="125" swimtime="00:01:09.17" />
                    <SPLIT distance="150" swimtime="00:01:25.58" />
                    <SPLIT distance="175" swimtime="00:01:39.87" />
                    <SPLIT distance="200" swimtime="00:01:52.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="4" lane="1" heat="1" heatid="10137" swimtime="00:04:00.45" reactiontime="+65" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:00:53.98" />
                    <SPLIT distance="125" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:25.52" />
                    <SPLIT distance="175" swimtime="00:01:41.18" />
                    <SPLIT distance="200" swimtime="00:01:57.12" />
                    <SPLIT distance="225" swimtime="00:02:12.91" />
                    <SPLIT distance="250" swimtime="00:02:29.93" />
                    <SPLIT distance="275" swimtime="00:02:47.30" />
                    <SPLIT distance="300" swimtime="00:03:04.53" />
                    <SPLIT distance="325" swimtime="00:03:19.09" />
                    <SPLIT distance="350" swimtime="00:03:32.88" />
                    <SPLIT distance="375" swimtime="00:03:46.84" />
                    <SPLIT distance="400" swimtime="00:04:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="7" lane="5" heat="2" heatid="20037" swimtime="00:04:04.32" reactiontime="+66" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                    <SPLIT distance="75" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:00:55.70" />
                    <SPLIT distance="125" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:27.56" />
                    <SPLIT distance="175" swimtime="00:01:43.36" />
                    <SPLIT distance="200" swimtime="00:01:58.63" />
                    <SPLIT distance="225" swimtime="00:02:15.37" />
                    <SPLIT distance="250" swimtime="00:02:32.58" />
                    <SPLIT distance="275" swimtime="00:02:49.99" />
                    <SPLIT distance="300" swimtime="00:03:07.45" />
                    <SPLIT distance="325" swimtime="00:03:22.12" />
                    <SPLIT distance="350" swimtime="00:03:36.13" />
                    <SPLIT distance="375" swimtime="00:03:50.37" />
                    <SPLIT distance="400" swimtime="00:04:04.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154844" lastname="CIAMPI" firstname="Matteo" gender="M" birthdate="1996-11-03">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.76" eventid="44" heat="5" lane="2">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:03:37.86" eventid="24" heat="5" lane="3">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="17" lane="2" heat="5" heatid="50044" swimtime="00:01:43.51" reactiontime="+70" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.47" />
                    <SPLIT distance="50" swimtime="00:00:24.26" />
                    <SPLIT distance="75" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:00:50.60" />
                    <SPLIT distance="125" swimtime="00:01:03.76" />
                    <SPLIT distance="150" swimtime="00:01:16.99" />
                    <SPLIT distance="175" swimtime="00:01:30.44" />
                    <SPLIT distance="200" swimtime="00:01:43.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="124" place="8" lane="5" heat="1" heatid="10124" swimtime="00:03:38.98" reactiontime="+70" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:25.03" />
                    <SPLIT distance="75" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:00:52.05" />
                    <SPLIT distance="125" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:19.66" />
                    <SPLIT distance="175" swimtime="00:01:33.71" />
                    <SPLIT distance="200" swimtime="00:01:47.60" />
                    <SPLIT distance="225" swimtime="00:02:01.72" />
                    <SPLIT distance="250" swimtime="00:02:15.83" />
                    <SPLIT distance="275" swimtime="00:02:29.82" />
                    <SPLIT distance="300" swimtime="00:02:43.91" />
                    <SPLIT distance="325" swimtime="00:02:57.97" />
                    <SPLIT distance="350" swimtime="00:03:12.00" />
                    <SPLIT distance="375" swimtime="00:03:25.82" />
                    <SPLIT distance="400" swimtime="00:03:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="2" lane="3" heat="5" heatid="50024" swimtime="00:03:37.73" reactiontime="+68" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:25.19" />
                    <SPLIT distance="75" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:00:52.37" />
                    <SPLIT distance="125" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:19.74" />
                    <SPLIT distance="175" swimtime="00:01:33.44" />
                    <SPLIT distance="200" swimtime="00:01:47.29" />
                    <SPLIT distance="225" swimtime="00:02:01.21" />
                    <SPLIT distance="250" swimtime="00:02:14.97" />
                    <SPLIT distance="275" swimtime="00:02:28.83" />
                    <SPLIT distance="300" swimtime="00:02:42.76" />
                    <SPLIT distance="325" swimtime="00:02:56.75" />
                    <SPLIT distance="350" swimtime="00:03:10.62" />
                    <SPLIT distance="375" swimtime="00:03:24.29" />
                    <SPLIT distance="400" swimtime="00:03:37.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149647" lastname="DEPLANO" firstname="Leonardo" gender="M" birthdate="1999-07-21">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.27" eventid="31" heat="9" lane="7">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="15" lane="7" heat="9" heatid="90031" swimtime="00:00:21.25" reactiontime="+68" points="853">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="12" lane="1" heat="1" heatid="10231" swimtime="00:00:21.12" reactiontime="+74" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.18" />
                    <SPLIT distance="50" swimtime="00:00:21.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119960" lastname="PANZIERA" firstname="Margherita" gender="F" birthdate="1995-08-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.51" eventid="2" heat="6" lane="7">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.05" eventid="45" heat="4" lane="5">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.22" eventid="18" heat="4" lane="6">
                  <MEETINFO date="2022-04-10" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="19" lane="7" heat="6" heatid="60002" swimtime="00:00:57.72" reactiontime="+57" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.71" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:00:57.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="5" lane="6" heat="1" heatid="10145" swimtime="00:02:02.18" reactiontime="+62" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.16" />
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="75" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:00:59.70" />
                    <SPLIT distance="125" swimtime="00:01:15.06" />
                    <SPLIT distance="150" swimtime="00:01:30.74" />
                    <SPLIT distance="175" swimtime="00:01:46.66" />
                    <SPLIT distance="200" swimtime="00:02:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="4" lane="5" heat="4" heatid="40045" swimtime="00:02:02.88" reactiontime="+62" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="75" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:00.23" />
                    <SPLIT distance="125" swimtime="00:01:15.83" />
                    <SPLIT distance="150" swimtime="00:01:31.58" />
                    <SPLIT distance="175" swimtime="00:01:47.47" />
                    <SPLIT distance="200" swimtime="00:02:02.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="26" lane="6" heat="4" heatid="40018" swimtime="00:00:27.30" reactiontime="+62" points="793">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="131052" lastname="SCALIA" firstname="Silvia" gender="F" birthdate="1995-07-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.78" eventid="2" heat="6" lane="6">
                  <MEETINFO date="2022-11-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:26.18" eventid="18" heat="5" lane="3">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="16" lane="6" heat="6" heatid="60002" swimtime="00:00:57.54" reactiontime="+57" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                    <SPLIT distance="75" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:00:57.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="16" lane="8" heat="1" heatid="10202" swimtime="00:00:58.02" reactiontime="+56" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                    <SPLIT distance="75" swimtime="00:00:42.70" />
                    <SPLIT distance="100" swimtime="00:00:58.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="13" lane="3" heat="5" heatid="50018" swimtime="00:00:26.40" reactiontime="+59" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="13" lane="1" heat="2" heatid="20218" swimtime="00:00:26.39" reactiontime="+61" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:26.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165018" lastname="PILATO" firstname="Benedetta" gender="F" birthdate="2005-01-18">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.66" eventid="15" heat="6" lane="3">
                  <MEETINFO date="2022-11-10" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.50" eventid="40" heat="6" lane="5">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="13" lane="3" heat="6" heatid="60015" swimtime="00:01:05.21" reactiontime="+70" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="75" swimtime="00:00:47.61" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="15" lane="1" heat="2" heatid="20215" swimtime="00:01:05.46" reactiontime="+68" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.63" />
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                    <SPLIT distance="75" swimtime="00:00:47.21" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="7" lane="7" heat="1" heatid="10140" swimtime="00:00:29.48" reactiontime="+65" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="7" lane="5" heat="6" heatid="60040" swimtime="00:00:29.63" reactiontime="+68" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="6" lane="6" heat="2" heatid="20240" swimtime="00:00:29.42" reactiontime="+66" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124777" lastname="CUSINATO" firstname="Ilaria" gender="F" birthdate="1999-10-05">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.30" eventid="20" heat="4" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:04:29.37" eventid="36" heat="3" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="10" lane="3" heat="4" heatid="40020" swimtime="00:02:06.01" reactiontime="+70" points="855">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="75" swimtime="00:00:43.90" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="125" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:32.40" />
                    <SPLIT distance="175" swimtime="00:01:49.12" />
                    <SPLIT distance="200" swimtime="00:02:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="7" lane="7" heat="1" heatid="10136" swimtime="00:04:32.68" reactiontime="+69" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="75" swimtime="00:00:45.87" />
                    <SPLIT distance="100" swimtime="00:01:02.74" />
                    <SPLIT distance="125" swimtime="00:01:20.60" />
                    <SPLIT distance="150" swimtime="00:01:37.76" />
                    <SPLIT distance="175" swimtime="00:01:55.04" />
                    <SPLIT distance="200" swimtime="00:02:11.91" />
                    <SPLIT distance="225" swimtime="00:02:31.28" />
                    <SPLIT distance="250" swimtime="00:02:50.88" />
                    <SPLIT distance="275" swimtime="00:03:10.38" />
                    <SPLIT distance="300" swimtime="00:03:30.09" />
                    <SPLIT distance="325" swimtime="00:03:46.52" />
                    <SPLIT distance="350" swimtime="00:04:01.99" />
                    <SPLIT distance="375" swimtime="00:04:17.67" />
                    <SPLIT distance="400" swimtime="00:04:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="6" lane="5" heat="3" heatid="30036" swimtime="00:04:32.94" reactiontime="+69" points="853">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                    <SPLIT distance="75" swimtime="00:00:45.35" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="125" swimtime="00:01:19.33" />
                    <SPLIT distance="150" swimtime="00:01:36.18" />
                    <SPLIT distance="175" swimtime="00:01:53.09" />
                    <SPLIT distance="200" swimtime="00:02:09.81" />
                    <SPLIT distance="225" swimtime="00:02:29.31" />
                    <SPLIT distance="250" swimtime="00:02:48.88" />
                    <SPLIT distance="275" swimtime="00:03:08.48" />
                    <SPLIT distance="300" swimtime="00:03:28.43" />
                    <SPLIT distance="325" swimtime="00:03:45.04" />
                    <SPLIT distance="350" swimtime="00:04:01.08" />
                    <SPLIT distance="375" swimtime="00:04:17.28" />
                    <SPLIT distance="400" swimtime="00:04:32.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124776" lastname="FRANCESCHI" firstname="Sara" gender="F" birthdate="1999-02-01">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.38" eventid="6" heat="4" lane="6">
                  <MEETINFO date="2022-11-10" />
                </ENTRY>
                <ENTRY entrytime="00:04:30.47" eventid="36" heat="4" lane="6">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="106" place="8" lane="8" heat="1" heatid="10106" swimtime="00:02:09.76" reactiontime="+72" points="828">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                    <SPLIT distance="75" swimtime="00:00:44.55" />
                    <SPLIT distance="100" swimtime="00:01:00.89" />
                    <SPLIT distance="125" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:01:38.21" />
                    <SPLIT distance="175" swimtime="00:01:54.59" />
                    <SPLIT distance="200" swimtime="00:02:09.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="8" lane="6" heat="4" heatid="40006" swimtime="00:02:07.25" reactiontime="+73" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="75" swimtime="00:00:44.57" />
                    <SPLIT distance="100" swimtime="00:00:59.88" />
                    <SPLIT distance="125" swimtime="00:01:17.87" />
                    <SPLIT distance="150" swimtime="00:01:36.27" />
                    <SPLIT distance="175" swimtime="00:01:52.51" />
                    <SPLIT distance="200" swimtime="00:02:07.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="2" lane="5" heat="1" heatid="10136" swimtime="00:04:28.58" reactiontime="+71" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.06" />
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="75" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:02.76" />
                    <SPLIT distance="125" swimtime="00:01:20.46" />
                    <SPLIT distance="150" swimtime="00:01:37.41" />
                    <SPLIT distance="175" swimtime="00:01:54.49" />
                    <SPLIT distance="200" swimtime="00:02:11.05" />
                    <SPLIT distance="225" swimtime="00:02:29.88" />
                    <SPLIT distance="250" swimtime="00:02:48.95" />
                    <SPLIT distance="275" swimtime="00:03:07.97" />
                    <SPLIT distance="300" swimtime="00:03:27.00" />
                    <SPLIT distance="325" swimtime="00:03:43.10" />
                    <SPLIT distance="350" swimtime="00:03:58.40" />
                    <SPLIT distance="375" swimtime="00:04:13.70" />
                    <SPLIT distance="400" swimtime="00:04:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="2" lane="6" heat="4" heatid="40036" swimtime="00:04:31.01" reactiontime="+73" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="75" swimtime="00:00:46.36" />
                    <SPLIT distance="100" swimtime="00:01:03.48" />
                    <SPLIT distance="125" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:01:37.86" />
                    <SPLIT distance="175" swimtime="00:01:54.84" />
                    <SPLIT distance="200" swimtime="00:02:12.14" />
                    <SPLIT distance="225" swimtime="00:02:30.35" />
                    <SPLIT distance="250" swimtime="00:02:49.32" />
                    <SPLIT distance="275" swimtime="00:03:08.41" />
                    <SPLIT distance="300" swimtime="00:03:27.76" />
                    <SPLIT distance="325" swimtime="00:03:44.28" />
                    <SPLIT distance="350" swimtime="00:04:00.20" />
                    <SPLIT distance="375" swimtime="00:04:16.04" />
                    <SPLIT distance="400" swimtime="00:04:31.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154343" lastname="COCCONCELLI" firstname="Costanza" gender="F" birthdate="2002-01-26">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.12" eventid="6" heat="4" lane="3">
                  <MEETINFO date="2022-11-10" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:58.45" eventid="22" heat="2" lane="5">
                  <MEETINFO date="2021-09-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="17" lane="3" heat="4" heatid="40006" swimtime="00:02:09.71" reactiontime="+65" points="829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:44.99" />
                    <SPLIT distance="100" swimtime="00:01:00.78" />
                    <SPLIT distance="125" swimtime="00:01:20.02" />
                    <SPLIT distance="150" swimtime="00:01:38.87" />
                    <SPLIT distance="175" swimtime="00:01:55.03" />
                    <SPLIT distance="200" swimtime="00:02:09.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="5" lane="5" heat="2" heatid="20022" swimtime="00:00:59.19" reactiontime="+63" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                    <SPLIT distance="75" swimtime="00:00:44.84" />
                    <SPLIT distance="100" swimtime="00:00:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="10" lane="3" heat="2" heatid="20222" swimtime="00:00:59.34" reactiontime="+63" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:00:59.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101725" lastname="DI PIETRO" firstname="Silvia" gender="F" birthdate="1993-04-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.03" eventid="4" heat="6" lane="3">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.94" eventid="30" heat="8" lane="6">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="8" lane="3" heat="6" heatid="60004" swimtime="00:00:25.32" reactiontime="+66" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="13" lane="2" heat="2" heatid="20204" swimtime="00:00:25.42" reactiontime="+67" points="882">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.81" />
                    <SPLIT distance="50" swimtime="00:00:25.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="-1" lane="6" heat="8" heatid="80030" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="190103" lastname="CONTE BONIN" firstname="Paolo" gender="M" birthdate="2002-02-09" />
            <ATHLETE athleteid="156605" lastname="FRIGO" firstname="Manuel" gender="M" birthdate="1997-02-18" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Italy">
              <RESULTS>
                <RESULT eventid="109" place="1" lane="4" heat="1" swimtime="00:03:02.75" reactiontime="+71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.45" />
                    <SPLIT distance="50" swimtime="00:00:22.06" />
                    <SPLIT distance="75" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:00:46.15" />
                    <SPLIT distance="125" swimtime="00:00:56.32" />
                    <SPLIT distance="150" swimtime="00:01:08.05" />
                    <SPLIT distance="175" swimtime="00:01:20.05" />
                    <SPLIT distance="200" swimtime="00:01:32.08" />
                    <SPLIT distance="225" swimtime="00:01:41.92" />
                    <SPLIT distance="250" swimtime="00:01:53.41" />
                    <SPLIT distance="275" swimtime="00:02:05.59" />
                    <SPLIT distance="300" swimtime="00:02:17.62" />
                    <SPLIT distance="325" swimtime="00:02:27.40" />
                    <SPLIT distance="350" swimtime="00:02:38.95" />
                    <SPLIT distance="375" swimtime="00:02:50.75" />
                    <SPLIT distance="400" swimtime="00:03:02.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124771" reactiontime="+71" />
                    <RELAYPOSITION number="2" athleteid="190103" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="149647" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="149646" reactiontime="+18" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="1" lane="4" heat="2" swimtime="00:03:04.46" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.42" />
                    <SPLIT distance="50" swimtime="00:00:22.03" />
                    <SPLIT distance="75" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:00:46.08" />
                    <SPLIT distance="125" swimtime="00:00:56.13" />
                    <SPLIT distance="150" swimtime="00:01:08.05" />
                    <SPLIT distance="175" swimtime="00:01:20.30" />
                    <SPLIT distance="200" swimtime="00:01:32.27" />
                    <SPLIT distance="225" swimtime="00:01:42.55" />
                    <SPLIT distance="250" swimtime="00:01:54.43" />
                    <SPLIT distance="275" swimtime="00:02:06.69" />
                    <SPLIT distance="300" swimtime="00:02:18.78" />
                    <SPLIT distance="325" swimtime="00:02:28.80" />
                    <SPLIT distance="350" swimtime="00:02:40.53" />
                    <SPLIT distance="375" swimtime="00:02:52.40" />
                    <SPLIT distance="400" swimtime="00:03:04.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124771" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="149647" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="156605" reactiontime="+30" />
                    <RELAYPOSITION number="4" athleteid="190103" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Italy">
              <RESULTS>
                <RESULT eventid="148" place="3" lane="3" heat="1" swimtime="00:03:19.06" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:23.89" />
                    <SPLIT distance="75" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:00:49.48" />
                    <SPLIT distance="125" swimtime="00:01:01.02" />
                    <SPLIT distance="150" swimtime="00:01:15.19" />
                    <SPLIT distance="175" swimtime="00:01:29.83" />
                    <SPLIT distance="200" swimtime="00:01:45.00" />
                    <SPLIT distance="225" swimtime="00:01:54.84" />
                    <SPLIT distance="250" swimtime="00:02:07.21" />
                    <SPLIT distance="275" swimtime="00:02:20.21" />
                    <SPLIT distance="300" swimtime="00:02:33.50" />
                    <SPLIT distance="325" swimtime="00:02:43.56" />
                    <SPLIT distance="350" swimtime="00:02:54.91" />
                    <SPLIT distance="375" swimtime="00:03:06.69" />
                    <SPLIT distance="400" swimtime="00:03:19.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154842" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="124772" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="102367" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="124771" reactiontime="+56" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="3" lane="4" heat="2" swimtime="00:03:23.81" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                    <SPLIT distance="50" swimtime="00:00:23.87" />
                    <SPLIT distance="75" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:00:49.59" />
                    <SPLIT distance="125" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:16.53" />
                    <SPLIT distance="175" swimtime="00:01:31.69" />
                    <SPLIT distance="200" swimtime="00:01:47.42" />
                    <SPLIT distance="225" swimtime="00:01:57.97" />
                    <SPLIT distance="250" swimtime="00:02:10.68" />
                    <SPLIT distance="275" swimtime="00:02:24.04" />
                    <SPLIT distance="300" swimtime="00:02:37.66" />
                    <SPLIT distance="325" swimtime="00:02:47.69" />
                    <SPLIT distance="350" swimtime="00:02:59.55" />
                    <SPLIT distance="375" swimtime="00:03:11.74" />
                    <SPLIT distance="400" swimtime="00:03:23.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="149646" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="198800" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="149648" reactiontime="+42" />
                    <RELAYPOSITION number="4" athleteid="190103" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Italy">
              <RESULTS>
                <RESULT eventid="132" place="3" lane="3" heat="1" swimtime="00:06:49.63" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.36" />
                    <SPLIT distance="50" swimtime="00:00:23.91" />
                    <SPLIT distance="75" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:00:50.04" />
                    <SPLIT distance="125" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:16.33" />
                    <SPLIT distance="175" swimtime="00:01:29.68" />
                    <SPLIT distance="200" swimtime="00:01:42.68" />
                    <SPLIT distance="225" swimtime="00:01:53.47" />
                    <SPLIT distance="250" swimtime="00:02:06.18" />
                    <SPLIT distance="275" swimtime="00:02:19.04" />
                    <SPLIT distance="300" swimtime="00:02:32.24" />
                    <SPLIT distance="325" swimtime="00:02:45.37" />
                    <SPLIT distance="350" swimtime="00:02:58.77" />
                    <SPLIT distance="375" swimtime="00:03:12.24" />
                    <SPLIT distance="400" swimtime="00:03:25.29" />
                    <SPLIT distance="425" swimtime="00:03:36.03" />
                    <SPLIT distance="450" swimtime="00:03:48.37" />
                    <SPLIT distance="475" swimtime="00:04:01.23" />
                    <SPLIT distance="500" swimtime="00:04:14.31" />
                    <SPLIT distance="525" swimtime="00:04:27.47" />
                    <SPLIT distance="550" swimtime="00:04:40.97" />
                    <SPLIT distance="575" swimtime="00:04:54.58" />
                    <SPLIT distance="600" swimtime="00:05:08.05" />
                    <SPLIT distance="625" swimtime="00:05:18.43" />
                    <SPLIT distance="650" swimtime="00:05:31.02" />
                    <SPLIT distance="675" swimtime="00:05:43.77" />
                    <SPLIT distance="700" swimtime="00:05:56.71" />
                    <SPLIT distance="725" swimtime="00:06:09.79" />
                    <SPLIT distance="750" swimtime="00:06:22.96" />
                    <SPLIT distance="775" swimtime="00:06:36.34" />
                    <SPLIT distance="800" swimtime="00:06:49.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154844" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="149646" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="149648" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="190103" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="3" lane="5" heat="2" swimtime="00:06:54.54" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.51" />
                    <SPLIT distance="50" swimtime="00:00:24.29" />
                    <SPLIT distance="75" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:00:50.51" />
                    <SPLIT distance="125" swimtime="00:01:03.79" />
                    <SPLIT distance="150" swimtime="00:01:17.08" />
                    <SPLIT distance="175" swimtime="00:01:30.43" />
                    <SPLIT distance="200" swimtime="00:01:43.50" />
                    <SPLIT distance="225" swimtime="00:01:54.27" />
                    <SPLIT distance="250" swimtime="00:02:07.03" />
                    <SPLIT distance="275" swimtime="00:02:20.38" />
                    <SPLIT distance="300" swimtime="00:02:33.81" />
                    <SPLIT distance="325" swimtime="00:02:47.07" />
                    <SPLIT distance="350" swimtime="00:03:00.58" />
                    <SPLIT distance="375" swimtime="00:03:14.16" />
                    <SPLIT distance="400" swimtime="00:03:27.56" />
                    <SPLIT distance="425" swimtime="00:03:38.17" />
                    <SPLIT distance="450" swimtime="00:03:50.80" />
                    <SPLIT distance="475" swimtime="00:04:03.83" />
                    <SPLIT distance="500" swimtime="00:04:16.86" />
                    <SPLIT distance="525" swimtime="00:04:30.10" />
                    <SPLIT distance="550" swimtime="00:04:43.65" />
                    <SPLIT distance="575" swimtime="00:04:57.41" />
                    <SPLIT distance="600" swimtime="00:05:10.84" />
                    <SPLIT distance="625" swimtime="00:05:21.85" />
                    <SPLIT distance="650" swimtime="00:05:34.49" />
                    <SPLIT distance="675" swimtime="00:05:47.55" />
                    <SPLIT distance="700" swimtime="00:06:00.80" />
                    <SPLIT distance="725" swimtime="00:06:14.33" />
                    <SPLIT distance="750" swimtime="00:06:27.90" />
                    <SPLIT distance="775" swimtime="00:06:41.46" />
                    <SPLIT distance="800" swimtime="00:06:54.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154844" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="156605" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="190103" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="149648" reactiontime="+47" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Italy">
              <RESULTS>
                <RESULT eventid="126" place="2" lane="3" heat="1" swimtime="00:01:23.48" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:21.22" />
                    <SPLIT distance="75" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:00:41.81" />
                    <SPLIT distance="125" swimtime="00:00:51.49" />
                    <SPLIT distance="150" swimtime="00:01:02.48" />
                    <SPLIT distance="175" swimtime="00:01:12.24" />
                    <SPLIT distance="200" swimtime="00:01:23.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124771" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="149647" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="149646" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="156605" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="3" lane="4" heat="1" swimtime="00:01:24.13" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.19" />
                    <SPLIT distance="50" swimtime="00:00:21.26" />
                    <SPLIT distance="75" swimtime="00:00:31.08" />
                    <SPLIT distance="100" swimtime="00:00:42.05" />
                    <SPLIT distance="125" swimtime="00:00:51.97" />
                    <SPLIT distance="150" swimtime="00:01:03.12" />
                    <SPLIT distance="175" swimtime="00:01:12.91" />
                    <SPLIT distance="200" swimtime="00:01:24.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124771" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="149647" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="156605" reactiontime="+33" />
                    <RELAYPOSITION number="4" athleteid="190103" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Italy">
              <RESULTS>
                <RESULT eventid="27" place="-1" lane="5" heat="4" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Italy">
              <RESULTS>
                <RESULT eventid="47" place="9" lane="3" heat="2" swimtime="00:03:55.62" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.32" />
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                    <SPLIT distance="75" swimtime="00:00:42.37" />
                    <SPLIT distance="100" swimtime="00:00:57.64" />
                    <SPLIT distance="125" swimtime="00:01:12.07" />
                    <SPLIT distance="150" swimtime="00:01:29.06" />
                    <SPLIT distance="175" swimtime="00:01:46.55" />
                    <SPLIT distance="200" swimtime="00:02:04.41" />
                    <SPLIT distance="225" swimtime="00:02:16.60" />
                    <SPLIT distance="250" swimtime="00:02:31.48" />
                    <SPLIT distance="275" swimtime="00:02:46.75" />
                    <SPLIT distance="300" swimtime="00:03:02.35" />
                    <SPLIT distance="325" swimtime="00:03:14.41" />
                    <SPLIT distance="350" swimtime="00:03:28.06" />
                    <SPLIT distance="375" swimtime="00:03:41.96" />
                    <SPLIT distance="400" swimtime="00:03:55.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="131052" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="124776" reactiontime="+41" />
                    <RELAYPOSITION number="3" athleteid="124777" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="154343" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Italy">
              <RESULTS>
                <RESULT eventid="34" place="-1" lane="3" heat="1" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Italy">
              <RESULTS>
                <RESULT eventid="111" place="2" lane="7" heat="1" swimtime="00:01:36.01" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.10" />
                    <SPLIT distance="50" swimtime="00:00:22.59" />
                    <SPLIT distance="75" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:00:47.42" />
                    <SPLIT distance="125" swimtime="00:00:58.41" />
                    <SPLIT distance="150" swimtime="00:01:11.94" />
                    <SPLIT distance="175" swimtime="00:01:23.46" />
                    <SPLIT distance="200" swimtime="00:01:36.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154842" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="124772" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="101725" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="154343" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="6" lane="4" heat="3" swimtime="00:01:38.91" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:23.17" />
                    <SPLIT distance="75" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:00:49.63" />
                    <SPLIT distance="125" swimtime="00:01:00.85" />
                    <SPLIT distance="150" swimtime="00:01:14.62" />
                    <SPLIT distance="175" swimtime="00:01:26.35" />
                    <SPLIT distance="200" swimtime="00:01:38.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154842" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="198800" reactiontime="+37" />
                    <RELAYPOSITION number="3" athleteid="101725" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="154343" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Italy">
              <RESULTS>
                <RESULT eventid="135" place="1" lane="4" heat="1" swimtime="00:01:29.72" reactiontime="+52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.09" />
                    <SPLIT distance="50" swimtime="00:00:22.65" />
                    <SPLIT distance="75" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:00:47.60" />
                    <SPLIT distance="125" swimtime="00:00:57.31" />
                    <SPLIT distance="150" swimtime="00:01:09.20" />
                    <SPLIT distance="175" swimtime="00:01:18.80" />
                    <SPLIT distance="200" swimtime="00:01:29.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154842" reactiontime="+52" />
                    <RELAYPOSITION number="2" athleteid="124772" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="102367" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="149647" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="1" lane="4" heat="3" swimtime="00:01:32.31" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:23.61" />
                    <SPLIT distance="75" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:00:49.67" />
                    <SPLIT distance="125" swimtime="00:00:59.38" />
                    <SPLIT distance="150" swimtime="00:01:11.47" />
                    <SPLIT distance="175" swimtime="00:01:21.38" />
                    <SPLIT distance="200" swimtime="00:01:32.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154842" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="198800" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="149646" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="124771" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Jamaica" shortname="JAM" code="JAM" nation="JAM" type="NOC">
          <ATHLETES />
        </CLUB>
        <CLUB name="Japan" shortname="JPN" code="JPN" nation="JPN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="101144" lastname="IRIE" firstname="Ryosuke" gender="M" birthdate="1990-01-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.66" eventid="3" heat="5" lane="5">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.21" eventid="19" heat="6" lane="6">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="10" lane="5" heat="5" heatid="50003" swimtime="00:00:50.37" reactiontime="+54" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:24.09" />
                    <SPLIT distance="75" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:00:50.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="9" lane="7" heat="2" heatid="20203" swimtime="00:00:50.08" reactiontime="+54" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:00:50.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="16" lane="6" heat="6" heatid="60019" swimtime="00:00:23.38" reactiontime="+53" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:23.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="14" lane="8" heat="1" heatid="10219" swimtime="00:00:23.49" reactiontime="+54" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:23.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214383" lastname="YANAGAWA" firstname="Daiki" gender="M" birthdate="2002-05-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.25" eventid="3" heat="4" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.94" eventid="46" heat="3" lane="6">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="19" lane="7" heat="4" heatid="40003" swimtime="00:00:50.99" reactiontime="+60" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                    <SPLIT distance="50" swimtime="00:00:24.94" />
                    <SPLIT distance="75" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:00:50.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="-1" lane="6" heat="3" heatid="30046" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129138" lastname="WATANABE" firstname="Ippei" gender="M" birthdate="1997-03-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.88" eventid="16" heat="6" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.70" eventid="29" heat="4" lane="4">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="6" lane="3" heat="6" heatid="60016" swimtime="00:00:57.11" reactiontime="+65" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                    <SPLIT distance="75" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="9" lane="3" heat="1" heatid="10216" swimtime="00:00:57.27" reactiontime="+64" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="75" swimtime="00:00:41.92" />
                    <SPLIT distance="100" swimtime="00:00:57.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="129" place="4" lane="3" heat="1" heatid="10129" swimtime="00:02:02.53" reactiontime="+66" points="943">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.52" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:43.33" />
                    <SPLIT distance="100" swimtime="00:00:58.86" />
                    <SPLIT distance="125" swimtime="00:01:14.68" />
                    <SPLIT distance="150" swimtime="00:01:30.47" />
                    <SPLIT distance="175" swimtime="00:01:46.39" />
                    <SPLIT distance="200" swimtime="00:02:02.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="3" lane="4" heat="4" heatid="40029" swimtime="00:02:03.64" reactiontime="+67" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.64" />
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="75" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:00:59.37" />
                    <SPLIT distance="125" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:31.46" />
                    <SPLIT distance="175" swimtime="00:01:47.75" />
                    <SPLIT distance="200" swimtime="00:02:03.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191038" lastname="HINOMOTO" firstname="Yuya" gender="M" birthdate="1997-02-14">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.77" eventid="16" heat="6" lane="4">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:26.09" eventid="41" heat="7" lane="5">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="8" lane="7" heat="1" heatid="10116" swimtime="00:00:57.29" reactiontime="+62" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="75" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:00:57.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="2" lane="4" heat="6" heatid="60016" swimtime="00:00:56.62" reactiontime="+65" points="930">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.08" />
                    <SPLIT distance="50" swimtime="00:00:26.39" />
                    <SPLIT distance="75" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="6" lane="4" heat="1" heatid="10216" swimtime="00:00:56.77" reactiontime="+61" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.14" />
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                    <SPLIT distance="75" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:00:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="6" lane="5" heat="7" heatid="70041" swimtime="00:00:26.15" reactiontime="+59" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="9" lane="3" heat="1" heatid="10241" swimtime="00:00:26.13" reactiontime="+61" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149684" lastname="SAKAMOTO" firstname="Yuya" gender="M" birthdate="1999-10-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.93" eventid="39" heat="6" lane="2">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="9" lane="2" heat="6" heatid="60039" swimtime="00:00:50.09" reactiontime="+64" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.62" />
                    <SPLIT distance="50" swimtime="00:00:23.57" />
                    <SPLIT distance="75" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:00:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="10" lane="2" heat="2" heatid="20239" swimtime="00:00:50.16" reactiontime="+64" points="864">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.55" />
                    <SPLIT distance="75" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:00:50.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214386" lastname="TANAKA" firstname="Yuya" gender="M" birthdate="1998-08-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.72" eventid="39" heat="7" lane="6">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.52" eventid="5" heat="8" lane="2">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="10" lane="6" heat="7" heatid="70039" swimtime="00:00:50.22" reactiontime="+61" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:23.09" />
                    <SPLIT distance="75" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:00:50.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="11" lane="2" heat="1" heatid="10239" swimtime="00:00:50.21" reactiontime="+60" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.59" />
                    <SPLIT distance="50" swimtime="00:00:23.15" />
                    <SPLIT distance="75" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:00:50.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="18" lane="2" heat="8" heatid="80005" swimtime="00:00:22.54" reactiontime="+59" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:22.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108761" lastname="NAKAMURA" firstname="Katsumi" gender="M" birthdate="1994-02-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.49" eventid="14" heat="9" lane="3">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="37" lane="3" heat="9" heatid="90014" swimtime="00:00:47.79" reactiontime="+71" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.84" />
                    <SPLIT distance="50" swimtime="00:00:22.92" />
                    <SPLIT distance="75" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130459" lastname="MATSUMOTO" firstname="Katsuhiro" gender="M" birthdate="1997-02-28">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.84" eventid="14" heat="11" lane="7">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.67" eventid="44" heat="5" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:03:39.54" eventid="24" heat="4" lane="2">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="22" lane="7" heat="11" heatid="110014" swimtime="00:00:47.13" reactiontime="+64" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.67" />
                    <SPLIT distance="50" swimtime="00:00:22.66" />
                    <SPLIT distance="75" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:00:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="144" place="8" lane="5" heat="1" heatid="10144" swimtime="00:01:41.91" reactiontime="+65" points="927">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.01" />
                    <SPLIT distance="50" swimtime="00:00:23.32" />
                    <SPLIT distance="75" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:00:49.29" />
                    <SPLIT distance="125" swimtime="00:01:02.38" />
                    <SPLIT distance="150" swimtime="00:01:15.57" />
                    <SPLIT distance="175" swimtime="00:01:28.74" />
                    <SPLIT distance="200" swimtime="00:01:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="2" lane="5" heat="5" heatid="50044" swimtime="00:01:41.29" reactiontime="+65" points="944">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.06" />
                    <SPLIT distance="50" swimtime="00:00:23.46" />
                    <SPLIT distance="75" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:00:49.17" />
                    <SPLIT distance="125" swimtime="00:01:02.29" />
                    <SPLIT distance="150" swimtime="00:01:15.25" />
                    <SPLIT distance="175" swimtime="00:01:28.41" />
                    <SPLIT distance="200" swimtime="00:01:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="124" place="4" lane="3" heat="1" heatid="10124" swimtime="00:03:36.87" reactiontime="+65" points="937">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:24.39" />
                    <SPLIT distance="75" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:00:51.46" />
                    <SPLIT distance="125" swimtime="00:01:05.17" />
                    <SPLIT distance="150" swimtime="00:01:18.94" />
                    <SPLIT distance="175" swimtime="00:01:32.88" />
                    <SPLIT distance="200" swimtime="00:01:46.94" />
                    <SPLIT distance="225" swimtime="00:02:00.75" />
                    <SPLIT distance="250" swimtime="00:02:14.44" />
                    <SPLIT distance="275" swimtime="00:02:28.22" />
                    <SPLIT distance="300" swimtime="00:02:42.05" />
                    <SPLIT distance="325" swimtime="00:02:55.90" />
                    <SPLIT distance="350" swimtime="00:03:09.68" />
                    <SPLIT distance="375" swimtime="00:03:23.57" />
                    <SPLIT distance="400" swimtime="00:03:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="3" lane="2" heat="4" heatid="40024" swimtime="00:03:37.96" reactiontime="+65" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.51" />
                    <SPLIT distance="50" swimtime="00:00:24.73" />
                    <SPLIT distance="75" swimtime="00:00:38.26" />
                    <SPLIT distance="100" swimtime="00:00:51.88" />
                    <SPLIT distance="125" swimtime="00:01:05.56" />
                    <SPLIT distance="150" swimtime="00:01:19.35" />
                    <SPLIT distance="175" swimtime="00:01:33.24" />
                    <SPLIT distance="200" swimtime="00:01:47.22" />
                    <SPLIT distance="225" swimtime="00:02:01.22" />
                    <SPLIT distance="250" swimtime="00:02:15.37" />
                    <SPLIT distance="275" swimtime="00:02:29.48" />
                    <SPLIT distance="300" swimtime="00:02:43.72" />
                    <SPLIT distance="325" swimtime="00:02:57.49" />
                    <SPLIT distance="350" swimtime="00:03:11.16" />
                    <SPLIT distance="375" swimtime="00:03:24.67" />
                    <SPLIT distance="400" swimtime="00:03:37.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108755" lastname="TAKEDA" firstname="Shogo" gender="M" birthdate="1995-01-01">
              <ENTRIES>
                <ENTRY entrytime="00:14:29.92" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:03:40.05" eventid="24" heat="4" lane="7">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="00:07:41.04" eventid="42" heat="0" lane="-1">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="4" lane="6" heat="5" heatid="30110" swimtime="00:14:25.95" reactiontime="+70" points="935">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.45" />
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="75" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:00:54.45" />
                    <SPLIT distance="125" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:22.87" />
                    <SPLIT distance="175" swimtime="00:01:36.90" />
                    <SPLIT distance="200" swimtime="00:01:51.23" />
                    <SPLIT distance="225" swimtime="00:02:05.39" />
                    <SPLIT distance="250" swimtime="00:02:19.72" />
                    <SPLIT distance="275" swimtime="00:02:34.16" />
                    <SPLIT distance="300" swimtime="00:02:48.59" />
                    <SPLIT distance="325" swimtime="00:03:03.12" />
                    <SPLIT distance="350" swimtime="00:03:17.59" />
                    <SPLIT distance="375" swimtime="00:03:31.99" />
                    <SPLIT distance="400" swimtime="00:03:46.37" />
                    <SPLIT distance="425" swimtime="00:04:00.89" />
                    <SPLIT distance="450" swimtime="00:04:15.25" />
                    <SPLIT distance="475" swimtime="00:04:29.70" />
                    <SPLIT distance="500" swimtime="00:04:44.23" />
                    <SPLIT distance="525" swimtime="00:04:58.71" />
                    <SPLIT distance="550" swimtime="00:05:13.10" />
                    <SPLIT distance="575" swimtime="00:05:27.54" />
                    <SPLIT distance="600" swimtime="00:05:42.17" />
                    <SPLIT distance="625" swimtime="00:05:56.60" />
                    <SPLIT distance="650" swimtime="00:06:11.11" />
                    <SPLIT distance="675" swimtime="00:06:25.65" />
                    <SPLIT distance="700" swimtime="00:06:40.13" />
                    <SPLIT distance="725" swimtime="00:06:54.80" />
                    <SPLIT distance="750" swimtime="00:07:09.37" />
                    <SPLIT distance="775" swimtime="00:07:24.00" />
                    <SPLIT distance="800" swimtime="00:07:38.74" />
                    <SPLIT distance="825" swimtime="00:07:53.18" />
                    <SPLIT distance="850" swimtime="00:08:07.81" />
                    <SPLIT distance="875" swimtime="00:08:22.58" />
                    <SPLIT distance="900" swimtime="00:08:37.30" />
                    <SPLIT distance="925" swimtime="00:08:51.72" />
                    <SPLIT distance="950" swimtime="00:09:06.58" />
                    <SPLIT distance="975" swimtime="00:09:21.24" />
                    <SPLIT distance="1000" swimtime="00:09:36.06" />
                    <SPLIT distance="1025" swimtime="00:09:50.71" />
                    <SPLIT distance="1050" swimtime="00:10:05.41" />
                    <SPLIT distance="1075" swimtime="00:10:20.15" />
                    <SPLIT distance="1100" swimtime="00:10:34.94" />
                    <SPLIT distance="1125" swimtime="00:10:49.57" />
                    <SPLIT distance="1150" swimtime="00:11:04.23" />
                    <SPLIT distance="1175" swimtime="00:11:18.83" />
                    <SPLIT distance="1200" swimtime="00:11:33.44" />
                    <SPLIT distance="1225" swimtime="00:11:48.02" />
                    <SPLIT distance="1250" swimtime="00:12:02.83" />
                    <SPLIT distance="1275" swimtime="00:12:17.51" />
                    <SPLIT distance="1300" swimtime="00:12:32.08" />
                    <SPLIT distance="1325" swimtime="00:12:46.65" />
                    <SPLIT distance="1350" swimtime="00:13:01.25" />
                    <SPLIT distance="1375" swimtime="00:13:15.70" />
                    <SPLIT distance="1400" swimtime="00:13:30.12" />
                    <SPLIT distance="1425" swimtime="00:13:44.53" />
                    <SPLIT distance="1450" swimtime="00:13:58.87" />
                    <SPLIT distance="1475" swimtime="00:14:12.75" />
                    <SPLIT distance="1500" swimtime="00:14:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="14" lane="7" heat="4" heatid="40024" swimtime="00:03:42.16" reactiontime="+67" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:25.62" />
                    <SPLIT distance="75" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:00:53.27" />
                    <SPLIT distance="125" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:21.41" />
                    <SPLIT distance="175" swimtime="00:01:35.38" />
                    <SPLIT distance="200" swimtime="00:01:49.58" />
                    <SPLIT distance="225" swimtime="00:02:03.54" />
                    <SPLIT distance="250" swimtime="00:02:17.81" />
                    <SPLIT distance="275" swimtime="00:02:31.92" />
                    <SPLIT distance="300" swimtime="00:02:46.27" />
                    <SPLIT distance="325" swimtime="00:03:00.35" />
                    <SPLIT distance="350" swimtime="00:03:14.38" />
                    <SPLIT distance="375" swimtime="00:03:28.55" />
                    <SPLIT distance="400" swimtime="00:03:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="4" lane="8" heat="5" heatid="30142" swimtime="00:07:33.78" reactiontime="+74" points="933">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:26.19" />
                    <SPLIT distance="75" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:00:54.73" />
                    <SPLIT distance="125" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:23.60" />
                    <SPLIT distance="175" swimtime="00:01:37.80" />
                    <SPLIT distance="200" swimtime="00:01:52.21" />
                    <SPLIT distance="225" swimtime="00:02:06.48" />
                    <SPLIT distance="250" swimtime="00:02:20.82" />
                    <SPLIT distance="275" swimtime="00:02:35.17" />
                    <SPLIT distance="300" swimtime="00:02:49.63" />
                    <SPLIT distance="325" swimtime="00:03:04.01" />
                    <SPLIT distance="350" swimtime="00:03:18.50" />
                    <SPLIT distance="375" swimtime="00:03:32.78" />
                    <SPLIT distance="400" swimtime="00:03:47.18" />
                    <SPLIT distance="425" swimtime="00:04:01.49" />
                    <SPLIT distance="450" swimtime="00:04:16.00" />
                    <SPLIT distance="475" swimtime="00:04:30.35" />
                    <SPLIT distance="500" swimtime="00:04:44.85" />
                    <SPLIT distance="525" swimtime="00:04:59.08" />
                    <SPLIT distance="550" swimtime="00:05:13.47" />
                    <SPLIT distance="575" swimtime="00:05:28.01" />
                    <SPLIT distance="600" swimtime="00:05:42.44" />
                    <SPLIT distance="625" swimtime="00:05:56.81" />
                    <SPLIT distance="650" swimtime="00:06:11.03" />
                    <SPLIT distance="675" swimtime="00:06:25.27" />
                    <SPLIT distance="700" swimtime="00:06:39.48" />
                    <SPLIT distance="725" swimtime="00:06:53.53" />
                    <SPLIT distance="750" swimtime="00:07:07.55" />
                    <SPLIT distance="775" swimtime="00:07:21.07" />
                    <SPLIT distance="800" swimtime="00:07:33.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214382" lastname="OZAKI" firstname="Kenta" gender="M" birthdate="1999-12-20">
              <ENTRIES>
                <ENTRY entrytime="00:14:45.13" eventid="10" heat="2" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="13" lane="5" heat="2" heatid="20010" swimtime="00:14:58.30" reactiontime="+69" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.48" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="75" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:00:55.25" />
                    <SPLIT distance="125" swimtime="00:01:09.83" />
                    <SPLIT distance="150" swimtime="00:01:24.52" />
                    <SPLIT distance="175" swimtime="00:01:39.24" />
                    <SPLIT distance="200" swimtime="00:01:53.95" />
                    <SPLIT distance="225" swimtime="00:02:08.60" />
                    <SPLIT distance="250" swimtime="00:02:23.39" />
                    <SPLIT distance="275" swimtime="00:02:38.30" />
                    <SPLIT distance="300" swimtime="00:02:53.19" />
                    <SPLIT distance="325" swimtime="00:03:08.10" />
                    <SPLIT distance="350" swimtime="00:03:23.07" />
                    <SPLIT distance="375" swimtime="00:03:37.92" />
                    <SPLIT distance="400" swimtime="00:03:52.82" />
                    <SPLIT distance="425" swimtime="00:04:07.73" />
                    <SPLIT distance="450" swimtime="00:04:22.80" />
                    <SPLIT distance="475" swimtime="00:04:37.77" />
                    <SPLIT distance="500" swimtime="00:04:52.74" />
                    <SPLIT distance="525" swimtime="00:05:07.79" />
                    <SPLIT distance="550" swimtime="00:05:22.79" />
                    <SPLIT distance="575" swimtime="00:05:37.71" />
                    <SPLIT distance="600" swimtime="00:05:52.86" />
                    <SPLIT distance="625" swimtime="00:06:07.89" />
                    <SPLIT distance="650" swimtime="00:06:22.95" />
                    <SPLIT distance="675" swimtime="00:06:38.01" />
                    <SPLIT distance="700" swimtime="00:06:53.15" />
                    <SPLIT distance="725" swimtime="00:07:08.27" />
                    <SPLIT distance="750" swimtime="00:07:23.41" />
                    <SPLIT distance="775" swimtime="00:07:38.40" />
                    <SPLIT distance="800" swimtime="00:07:53.51" />
                    <SPLIT distance="825" swimtime="00:08:08.53" />
                    <SPLIT distance="850" swimtime="00:08:23.81" />
                    <SPLIT distance="875" swimtime="00:08:38.83" />
                    <SPLIT distance="900" swimtime="00:08:54.08" />
                    <SPLIT distance="925" swimtime="00:09:09.05" />
                    <SPLIT distance="950" swimtime="00:09:24.46" />
                    <SPLIT distance="975" swimtime="00:09:39.72" />
                    <SPLIT distance="1000" swimtime="00:09:54.79" />
                    <SPLIT distance="1025" swimtime="00:10:09.98" />
                    <SPLIT distance="1050" swimtime="00:10:25.28" />
                    <SPLIT distance="1075" swimtime="00:10:40.50" />
                    <SPLIT distance="1100" swimtime="00:10:55.87" />
                    <SPLIT distance="1125" swimtime="00:11:11.09" />
                    <SPLIT distance="1150" swimtime="00:11:26.62" />
                    <SPLIT distance="1175" swimtime="00:11:41.86" />
                    <SPLIT distance="1200" swimtime="00:11:57.36" />
                    <SPLIT distance="1225" swimtime="00:12:12.72" />
                    <SPLIT distance="1250" swimtime="00:12:28.49" />
                    <SPLIT distance="1275" swimtime="00:12:43.80" />
                    <SPLIT distance="1300" swimtime="00:12:59.29" />
                    <SPLIT distance="1325" swimtime="00:13:14.53" />
                    <SPLIT distance="1350" swimtime="00:13:30.33" />
                    <SPLIT distance="1375" swimtime="00:13:45.56" />
                    <SPLIT distance="1400" swimtime="00:14:00.68" />
                    <SPLIT distance="1425" swimtime="00:14:15.27" />
                    <SPLIT distance="1450" swimtime="00:14:30.34" />
                    <SPLIT distance="1475" swimtime="00:14:44.56" />
                    <SPLIT distance="1500" swimtime="00:14:58.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214385" lastname="NAITO" firstname="Ryota" gender="M" birthdate="1997-10-30">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.93" eventid="46" heat="2" lane="5">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="146" place="8" lane="1" heat="1" heatid="10146" swimtime="00:01:51.67" reactiontime="+60" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:00:53.45" />
                    <SPLIT distance="125" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:22.26" />
                    <SPLIT distance="175" swimtime="00:01:37.15" />
                    <SPLIT distance="200" swimtime="00:01:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="7" lane="5" heat="2" heatid="20046" swimtime="00:01:50.78" reactiontime="+59" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                    <SPLIT distance="75" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:00:53.27" />
                    <SPLIT distance="125" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:21.74" />
                    <SPLIT distance="175" swimtime="00:01:36.49" />
                    <SPLIT distance="200" swimtime="00:01:50.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100478" lastname="SETO" firstname="Daiya" gender="M" birthdate="1994-05-24">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.49" eventid="29" heat="5" lane="4">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:01:49.41" eventid="21" heat="3" lane="4">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.66" eventid="7" heat="4" lane="4">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:03:56.26" eventid="37" heat="3" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="129" place="1" lane="4" heat="1" heatid="10129" swimtime="00:02:00.35" reactiontime="+60" points="995">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.50" />
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                    <SPLIT distance="75" swimtime="00:00:42.93" />
                    <SPLIT distance="100" swimtime="00:00:58.44" />
                    <SPLIT distance="125" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:29.42" />
                    <SPLIT distance="175" swimtime="00:01:44.83" />
                    <SPLIT distance="200" swimtime="00:02:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="1" lane="4" heat="5" heatid="50029" swimtime="00:02:02.43" reactiontime="+61" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                    <SPLIT distance="75" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:00:59.35" />
                    <SPLIT distance="125" swimtime="00:01:14.94" />
                    <SPLIT distance="150" swimtime="00:01:30.71" />
                    <SPLIT distance="175" swimtime="00:01:46.67" />
                    <SPLIT distance="200" swimtime="00:02:02.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="121" place="2" lane="3" heat="1" heatid="10121" swimtime="00:01:49.22" reactiontime="+61" points="973">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.96" />
                    <SPLIT distance="50" swimtime="00:00:24.41" />
                    <SPLIT distance="75" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:00:52.13" />
                    <SPLIT distance="125" swimtime="00:01:05.94" />
                    <SPLIT distance="150" swimtime="00:01:20.15" />
                    <SPLIT distance="175" swimtime="00:01:34.41" />
                    <SPLIT distance="200" swimtime="00:01:49.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="3" lane="4" heat="3" heatid="30021" swimtime="00:01:49.99" reactiontime="+63" points="953">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.15" />
                    <SPLIT distance="50" swimtime="00:00:24.73" />
                    <SPLIT distance="75" swimtime="00:00:38.95" />
                    <SPLIT distance="100" swimtime="00:00:53.01" />
                    <SPLIT distance="125" swimtime="00:01:07.01" />
                    <SPLIT distance="150" swimtime="00:01:21.11" />
                    <SPLIT distance="175" swimtime="00:01:35.51" />
                    <SPLIT distance="200" swimtime="00:01:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="107" place="5" lane="4" heat="1" heatid="10107" swimtime="00:01:51.39" reactiontime="+59" points="953">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.00" />
                    <SPLIT distance="50" swimtime="00:00:24.30" />
                    <SPLIT distance="75" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:00:52.28" />
                    <SPLIT distance="125" swimtime="00:01:08.03" />
                    <SPLIT distance="150" swimtime="00:01:24.05" />
                    <SPLIT distance="175" swimtime="00:01:38.21" />
                    <SPLIT distance="200" swimtime="00:01:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="1" lane="4" heat="4" heatid="40007" swimtime="00:01:51.76" reactiontime="+61" points="943">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.05" />
                    <SPLIT distance="50" swimtime="00:00:24.20" />
                    <SPLIT distance="75" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                    <SPLIT distance="125" swimtime="00:01:08.34" />
                    <SPLIT distance="150" swimtime="00:01:24.33" />
                    <SPLIT distance="175" swimtime="00:01:38.50" />
                    <SPLIT distance="200" swimtime="00:01:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="1" lane="4" heat="1" heatid="10137" swimtime="00:03:55.75" reactiontime="+62" points="988">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.18" />
                    <SPLIT distance="50" swimtime="00:00:25.00" />
                    <SPLIT distance="75" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:00:53.69" />
                    <SPLIT distance="125" swimtime="00:01:08.73" />
                    <SPLIT distance="150" swimtime="00:01:23.48" />
                    <SPLIT distance="175" swimtime="00:01:38.53" />
                    <SPLIT distance="200" swimtime="00:01:53.29" />
                    <SPLIT distance="225" swimtime="00:02:09.43" />
                    <SPLIT distance="250" swimtime="00:02:25.93" />
                    <SPLIT distance="275" swimtime="00:02:42.33" />
                    <SPLIT distance="300" swimtime="00:02:58.83" />
                    <SPLIT distance="325" swimtime="00:03:13.34" />
                    <SPLIT distance="350" swimtime="00:03:27.39" />
                    <SPLIT distance="375" swimtime="00:03:41.65" />
                    <SPLIT distance="400" swimtime="00:03:55.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="1" lane="4" heat="3" heatid="30037" swimtime="00:04:00.35" reactiontime="+61" points="932">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:25.01" />
                    <SPLIT distance="75" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:00:53.95" />
                    <SPLIT distance="125" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:24.01" />
                    <SPLIT distance="175" swimtime="00:01:39.40" />
                    <SPLIT distance="200" swimtime="00:01:54.49" />
                    <SPLIT distance="225" swimtime="00:02:11.26" />
                    <SPLIT distance="250" swimtime="00:02:27.96" />
                    <SPLIT distance="275" swimtime="00:02:44.94" />
                    <SPLIT distance="300" swimtime="00:03:02.12" />
                    <SPLIT distance="325" swimtime="00:03:17.05" />
                    <SPLIT distance="350" swimtime="00:03:31.52" />
                    <SPLIT distance="375" swimtime="00:03:46.19" />
                    <SPLIT distance="400" swimtime="00:04:00.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214387" lastname="MORIMOTO" firstname="Teppei" gender="M" birthdate="2002-04-07">
              <ENTRIES>
                <ENTRY entrytime="00:01:50.44" eventid="21" heat="4" lane="3">
                  <MEETINFO date="2021-12-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="121" place="6" lane="6" heat="1" heatid="10121" swimtime="00:01:50.70" reactiontime="+64" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:24.95" />
                    <SPLIT distance="75" swimtime="00:00:39.27" />
                    <SPLIT distance="100" swimtime="00:00:53.60" />
                    <SPLIT distance="125" swimtime="00:01:07.67" />
                    <SPLIT distance="150" swimtime="00:01:21.88" />
                    <SPLIT distance="175" swimtime="00:01:36.21" />
                    <SPLIT distance="200" swimtime="00:01:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="4" lane="3" heat="4" heatid="40021" swimtime="00:01:50.26" reactiontime="+62" points="946">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.26" />
                    <SPLIT distance="50" swimtime="00:00:24.94" />
                    <SPLIT distance="75" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:00:53.39" />
                    <SPLIT distance="125" swimtime="00:01:07.53" />
                    <SPLIT distance="150" swimtime="00:01:21.94" />
                    <SPLIT distance="175" swimtime="00:01:36.12" />
                    <SPLIT distance="200" swimtime="00:01:50.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214381" lastname="MANO" firstname="Hidenari" gender="M" birthdate="2000-07-06">
              <ENTRIES>
                <ENTRY entrytime="00:01:43.25" eventid="44" heat="4" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="19" lane="7" heat="4" heatid="40044" swimtime="00:01:44.20" reactiontime="+65" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:23.86" />
                    <SPLIT distance="75" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:00:50.09" />
                    <SPLIT distance="125" swimtime="00:01:03.40" />
                    <SPLIT distance="150" swimtime="00:01:16.95" />
                    <SPLIT distance="175" swimtime="00:01:30.69" />
                    <SPLIT distance="200" swimtime="00:01:44.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214388" lastname="OGATA" firstname="So" gender="M" birthdate="2003-04-28">
              <ENTRIES>
                <ENTRY entrytime="00:01:52.93" eventid="7" heat="3" lane="3">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:04:01.67" eventid="37" heat="2" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="107" place="8" lane="8" heat="1" heatid="10107" swimtime="00:01:53.40" reactiontime="+64" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.24" />
                    <SPLIT distance="50" swimtime="00:00:24.67" />
                    <SPLIT distance="75" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:00:53.03" />
                    <SPLIT distance="125" swimtime="00:01:09.31" />
                    <SPLIT distance="150" swimtime="00:01:26.02" />
                    <SPLIT distance="175" swimtime="00:01:40.47" />
                    <SPLIT distance="200" swimtime="00:01:53.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="8" lane="3" heat="3" heatid="30007" swimtime="00:01:53.00" reactiontime="+63" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                    <SPLIT distance="75" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:00:53.14" />
                    <SPLIT distance="125" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:25.79" />
                    <SPLIT distance="175" swimtime="00:01:39.99" />
                    <SPLIT distance="200" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="5" lane="7" heat="1" heatid="10137" swimtime="00:04:02.21" reactiontime="+66" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:25.80" />
                    <SPLIT distance="75" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:00:55.10" />
                    <SPLIT distance="125" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:26.18" />
                    <SPLIT distance="175" swimtime="00:01:41.48" />
                    <SPLIT distance="200" swimtime="00:01:56.22" />
                    <SPLIT distance="225" swimtime="00:02:13.11" />
                    <SPLIT distance="250" swimtime="00:02:30.28" />
                    <SPLIT distance="275" swimtime="00:02:47.61" />
                    <SPLIT distance="300" swimtime="00:03:04.98" />
                    <SPLIT distance="325" swimtime="00:03:20.33" />
                    <SPLIT distance="350" swimtime="00:03:34.76" />
                    <SPLIT distance="375" swimtime="00:03:48.94" />
                    <SPLIT distance="400" swimtime="00:04:02.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="6" lane="3" heat="2" heatid="20037" swimtime="00:04:03.29" reactiontime="+63" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.60" />
                    <SPLIT distance="50" swimtime="00:00:25.73" />
                    <SPLIT distance="75" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:00:54.95" />
                    <SPLIT distance="125" swimtime="00:01:11.02" />
                    <SPLIT distance="150" swimtime="00:01:26.09" />
                    <SPLIT distance="175" swimtime="00:01:41.36" />
                    <SPLIT distance="200" swimtime="00:01:56.10" />
                    <SPLIT distance="225" swimtime="00:02:12.83" />
                    <SPLIT distance="250" swimtime="00:02:29.92" />
                    <SPLIT distance="275" swimtime="00:02:47.48" />
                    <SPLIT distance="300" swimtime="00:03:04.75" />
                    <SPLIT distance="325" swimtime="00:03:20.24" />
                    <SPLIT distance="350" swimtime="00:03:34.71" />
                    <SPLIT distance="375" swimtime="00:03:49.19" />
                    <SPLIT distance="400" swimtime="00:04:03.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118529" lastname="KAWAMOTO" firstname="Takeshi" gender="M" birthdate="1995-02-19">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.11" eventid="19" heat="6" lane="3">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.28" eventid="5" heat="8" lane="3">
                  <MEETINFO date="2021-08-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="11" lane="3" heat="6" heatid="60019" swimtime="00:00:23.25" reactiontime="+54" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:23.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="12" lane="7" heat="1" heatid="10219" swimtime="00:00:23.19" reactiontime="+58" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:23.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="11" lane="3" heat="8" heatid="80005" swimtime="00:00:22.38" reactiontime="+59" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.37" />
                    <SPLIT distance="50" swimtime="00:00:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="15" lane="7" heat="2" heatid="20205" swimtime="00:00:22.50" reactiontime="+63" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.38" />
                    <SPLIT distance="50" swimtime="00:00:22.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157430" lastname="NIIYAMA" firstname="Masaki" gender="M" birthdate="1993-06-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.16" eventid="41" heat="8" lane="6">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="16" lane="6" heat="8" heatid="80041" swimtime="00:00:26.51" reactiontime="+62" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="341" place="17" lane="4" heat="1" heatid="10341" swimtime="00:00:26.50" reactiontime="+60" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:26.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130485" lastname="MATSUI" firstname="Kosuke" gender="M" birthdate="1994-03-28">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.16" eventid="31" heat="11" lane="6">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="12" lane="6" heat="11" heatid="110031" swimtime="00:00:21.17" reactiontime="+56" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.03" />
                    <SPLIT distance="50" swimtime="00:00:21.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="16" lane="7" heat="1" heatid="10231" swimtime="00:00:21.42" reactiontime="+59" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.11" />
                    <SPLIT distance="50" swimtime="00:00:21.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214380" lastname="KAWANE" firstname="Masahiro" gender="M" birthdate="1999-07-18">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.18" eventid="31" heat="11" lane="2">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="34" lane="2" heat="11" heatid="110031" swimtime="00:00:21.55" reactiontime="+61" points="818">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.41" />
                    <SPLIT distance="50" swimtime="00:00:21.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101276" lastname="AKASE" firstname="Sayaka" gender="F" birthdate="1994-08-25">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.04" eventid="2" heat="6" lane="1">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.72" eventid="45" heat="5" lane="2">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="14" lane="1" heat="6" heatid="60002" swimtime="00:00:57.51" reactiontime="+56" points="869">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.49" />
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="75" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="15" lane="8" heat="2" heatid="20202" swimtime="00:00:57.65" reactiontime="+56" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="75" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:00:57.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="15" lane="2" heat="5" heatid="50045" swimtime="00:02:05.13" reactiontime="+57" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.16" />
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="75" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:01.56" />
                    <SPLIT distance="125" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:01:33.46" />
                    <SPLIT distance="175" swimtime="00:01:49.40" />
                    <SPLIT distance="200" swimtime="00:02:05.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153984" lastname="SHIRAI" firstname="Rio" gender="F" birthdate="1999-09-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.91" eventid="2" heat="5" lane="6">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.85" eventid="13" heat="7" lane="2">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="18" lane="6" heat="5" heatid="50002" swimtime="00:00:57.71" reactiontime="+56" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="75" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:00:57.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="24" lane="2" heat="7" heatid="70013" swimtime="00:00:53.88" reactiontime="+70" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:26.06" />
                    <SPLIT distance="75" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:00:53.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130477" lastname="AOKI" firstname="Reona" gender="F" birthdate="1995-02-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.01" eventid="15" heat="6" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:29.59" eventid="40" heat="7" lane="3">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="6" lane="3" heat="1" heatid="10115" swimtime="00:01:04.30" reactiontime="+59" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.83" />
                    <SPLIT distance="50" swimtime="00:00:30.04" />
                    <SPLIT distance="75" swimtime="00:00:46.96" />
                    <SPLIT distance="100" swimtime="00:01:04.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="8" lane="5" heat="6" heatid="60015" swimtime="00:01:04.58" reactiontime="+65" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="75" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:04.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="3" lane="6" heat="1" heatid="10215" swimtime="00:01:04.13" reactiontime="+63" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.64" />
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="75" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="10" lane="3" heat="7" heatid="70040" swimtime="00:00:29.81" reactiontime="+63" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.85" />
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="12" lane="2" heat="1" heatid="10240" swimtime="00:00:30.01" reactiontime="+58" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214389" lastname="FUKASAWA" firstname="Mai" gender="F" birthdate="1998-10-15">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.00" eventid="15" heat="6" lane="2">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="7" lane="1" heat="1" heatid="10115" swimtime="00:01:04.48" reactiontime="+62" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.42" />
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="75" swimtime="00:00:47.35" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="7" lane="2" heat="6" heatid="60015" swimtime="00:01:04.57" reactiontime="+62" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="75" swimtime="00:00:47.58" />
                    <SPLIT distance="100" swimtime="00:01:04.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="7" lane="6" heat="2" heatid="20215" swimtime="00:01:04.45" reactiontime="+66" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.30" />
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="75" swimtime="00:00:47.48" />
                    <SPLIT distance="100" swimtime="00:01:04.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153983" lastname="SOMA" firstname="Ai" gender="F" birthdate="1997-09-15">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:56.68" eventid="38" heat="3" lane="3">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.07" eventid="4" heat="5" lane="3">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="138" place="5" lane="8" heat="1" heatid="10138" swimtime="00:00:56.27" reactiontime="+66" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="75" swimtime="00:00:40.83" />
                    <SPLIT distance="100" swimtime="00:00:56.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="7" lane="3" heat="3" heatid="30038" swimtime="00:00:56.72" reactiontime="+65" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                    <SPLIT distance="75" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:00:56.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="9" lane="6" heat="2" heatid="20238" swimtime="00:00:56.51" reactiontime="+68" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.08" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="75" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:00:56.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="8" lane="3" heat="5" heatid="50004" swimtime="00:00:25.32" reactiontime="+62" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                    <SPLIT distance="50" swimtime="00:00:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="10" lane="6" heat="1" heatid="10204" swimtime="00:00:25.36" reactiontime="+63" points="888">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214391" lastname="TSUDA" firstname="Moe" gender="F" birthdate="2000-12-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.71" eventid="38" heat="2" lane="3">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.26" eventid="4" heat="6" lane="6">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="12" lane="3" heat="2" heatid="20038" swimtime="00:00:57.22" reactiontime="+60" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="75" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:00:57.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="15" lane="7" heat="1" heatid="10238" swimtime="00:00:57.25" reactiontime="+63" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:26.98" />
                    <SPLIT distance="75" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:00:57.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="12" lane="6" heat="6" heatid="60004" swimtime="00:00:25.47" reactiontime="+61" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                    <SPLIT distance="50" swimtime="00:00:25.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="12" lane="7" heat="1" heatid="10204" swimtime="00:00:25.41" reactiontime="+62" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.67" />
                    <SPLIT distance="50" swimtime="00:00:25.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100703" lastname="IGARASHI" firstname="Chihiro" gender="F" birthdate="1995-05-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:52.84" eventid="13" heat="8" lane="2">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.34" eventid="43" heat="5" lane="2">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="17" lane="2" heat="8" heatid="80013" swimtime="00:00:53.38" reactiontime="+58" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.19" />
                    <SPLIT distance="50" swimtime="00:00:25.74" />
                    <SPLIT distance="75" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:00:53.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="14" lane="2" heat="5" heatid="50043" swimtime="00:01:56.22" reactiontime="+58" points="855">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                    <SPLIT distance="75" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:00:56.46" />
                    <SPLIT distance="125" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:26.59" />
                    <SPLIT distance="175" swimtime="00:01:41.75" />
                    <SPLIT distance="200" swimtime="00:01:56.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210159" lastname="YAMAMOTO" firstname="Chiaki" gender="F" birthdate="2007-03-08">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.66" eventid="45" heat="3" lane="6">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="18" lane="6" heat="3" heatid="30045" swimtime="00:02:06.10" reactiontime="+60" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="75" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="125" swimtime="00:01:17.58" />
                    <SPLIT distance="150" swimtime="00:01:33.95" />
                    <SPLIT distance="175" swimtime="00:01:50.51" />
                    <SPLIT distance="200" swimtime="00:02:06.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210164" lastname="KUSUDA" firstname="Yumeno" gender="F" birthdate="2005-10-25">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.36" eventid="28" heat="5" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="12" lane="7" heat="5" heatid="50028" swimtime="00:02:20.82" reactiontime="+72" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="75" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="125" swimtime="00:01:26.06" />
                    <SPLIT distance="150" swimtime="00:01:44.30" />
                    <SPLIT distance="175" swimtime="00:02:02.58" />
                    <SPLIT distance="200" swimtime="00:02:20.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214390" lastname="KATO" firstname="Kotomi" gender="F" birthdate="2006-01-05">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.89" eventid="28" heat="3" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="-1" lane="7" heat="3" heatid="30028" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214392" lastname="MITSUI" firstname="Airi" gender="F" birthdate="2004-06-12">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.35" eventid="20" heat="2" lane="4">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="120" place="6" lane="2" heat="1" heatid="10120" swimtime="00:02:05.40" reactiontime="+67" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                    <SPLIT distance="75" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:00.80" />
                    <SPLIT distance="125" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:01:32.82" />
                    <SPLIT distance="175" swimtime="00:01:48.94" />
                    <SPLIT distance="200" swimtime="00:02:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="5" lane="4" heat="2" heatid="20020" swimtime="00:02:05.27" reactiontime="+71" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="75" swimtime="00:00:45.30" />
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                    <SPLIT distance="125" swimtime="00:01:17.48" />
                    <SPLIT distance="150" swimtime="00:01:33.37" />
                    <SPLIT distance="175" swimtime="00:01:49.21" />
                    <SPLIT distance="200" swimtime="00:02:05.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214393" lastname="UCHIDA" firstname="Karin" gender="F" birthdate="2000-08-24">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.74" eventid="20" heat="4" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="120" place="7" lane="7" heat="1" heatid="10120" swimtime="00:02:05.51" reactiontime="+65" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="75" swimtime="00:00:44.18" />
                    <SPLIT distance="100" swimtime="00:01:00.49" />
                    <SPLIT distance="125" swimtime="00:01:16.53" />
                    <SPLIT distance="150" swimtime="00:01:32.89" />
                    <SPLIT distance="175" swimtime="00:01:49.20" />
                    <SPLIT distance="200" swimtime="00:02:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="6" lane="5" heat="4" heatid="40020" swimtime="00:02:05.38" reactiontime="+64" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.93" />
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                    <SPLIT distance="75" swimtime="00:00:44.30" />
                    <SPLIT distance="100" swimtime="00:01:00.39" />
                    <SPLIT distance="125" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:32.67" />
                    <SPLIT distance="175" swimtime="00:01:49.08" />
                    <SPLIT distance="200" swimtime="00:02:05.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130482" lastname="OHASHI" firstname="Yui" gender="F" birthdate="1995-10-18">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.86" eventid="6" heat="3" lane="4">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.05" eventid="22" heat="3" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="13" lane="4" heat="3" heatid="30006" swimtime="00:02:08.12" reactiontime="+67" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.74" />
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                    <SPLIT distance="75" swimtime="00:00:44.36" />
                    <SPLIT distance="100" swimtime="00:01:00.14" />
                    <SPLIT distance="125" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:01:37.43" />
                    <SPLIT distance="175" swimtime="00:01:53.53" />
                    <SPLIT distance="200" swimtime="00:02:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="10" lane="3" heat="3" heatid="30022" swimtime="00:00:59.49" reactiontime="+65" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                    <SPLIT distance="75" swimtime="00:00:44.94" />
                    <SPLIT distance="100" swimtime="00:00:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="11" lane="2" heat="1" heatid="10222" swimtime="00:00:59.45" reactiontime="+63" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                    <SPLIT distance="75" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:00:59.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214394" lastname="NAKASHIMA" firstname="Ao" gender="F" birthdate="2007-06-28">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.85" eventid="6" heat="5" lane="1">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="15" lane="1" heat="5" heatid="50006" swimtime="00:02:09.55" reactiontime="+65" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="75" swimtime="00:00:44.86" />
                    <SPLIT distance="100" swimtime="00:01:01.40" />
                    <SPLIT distance="125" swimtime="00:01:19.69" />
                    <SPLIT distance="150" swimtime="00:01:38.21" />
                    <SPLIT distance="175" swimtime="00:01:54.61" />
                    <SPLIT distance="200" swimtime="00:02:09.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149685" lastname="KOBORI" firstname="Waka" gender="F" birthdate="2000-08-10">
              <ENTRIES>
                <ENTRY entrytime="00:04:02.86" eventid="1" heat="4" lane="7">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="00:04:33.56" eventid="36" heat="3" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="101" place="7" lane="7" heat="1" heatid="10101" swimtime="00:04:02.14" reactiontime="+71" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:00:58.26" />
                    <SPLIT distance="125" swimtime="00:01:13.43" />
                    <SPLIT distance="150" swimtime="00:01:28.86" />
                    <SPLIT distance="175" swimtime="00:01:44.37" />
                    <SPLIT distance="200" swimtime="00:02:00.00" />
                    <SPLIT distance="225" swimtime="00:02:15.36" />
                    <SPLIT distance="250" swimtime="00:02:30.90" />
                    <SPLIT distance="275" swimtime="00:02:46.27" />
                    <SPLIT distance="300" swimtime="00:03:01.78" />
                    <SPLIT distance="325" swimtime="00:03:17.12" />
                    <SPLIT distance="350" swimtime="00:03:32.68" />
                    <SPLIT distance="375" swimtime="00:03:47.86" />
                    <SPLIT distance="400" swimtime="00:04:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="6" lane="7" heat="4" heatid="40001" swimtime="00:04:02.05" reactiontime="+70" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.41" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:00:58.37" />
                    <SPLIT distance="125" swimtime="00:01:13.54" />
                    <SPLIT distance="150" swimtime="00:01:28.94" />
                    <SPLIT distance="175" swimtime="00:01:44.07" />
                    <SPLIT distance="200" swimtime="00:01:59.56" />
                    <SPLIT distance="225" swimtime="00:02:14.66" />
                    <SPLIT distance="250" swimtime="00:02:30.14" />
                    <SPLIT distance="275" swimtime="00:02:45.35" />
                    <SPLIT distance="300" swimtime="00:03:01.00" />
                    <SPLIT distance="325" swimtime="00:03:16.44" />
                    <SPLIT distance="350" swimtime="00:03:32.06" />
                    <SPLIT distance="375" swimtime="00:03:47.20" />
                    <SPLIT distance="400" swimtime="00:04:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="3" lane="3" heat="1" heatid="10136" swimtime="00:04:29.03" reactiontime="+72" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="75" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="125" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                    <SPLIT distance="175" swimtime="00:01:54.61" />
                    <SPLIT distance="200" swimtime="00:02:11.38" />
                    <SPLIT distance="225" swimtime="00:02:30.63" />
                    <SPLIT distance="250" swimtime="00:02:49.93" />
                    <SPLIT distance="275" swimtime="00:03:09.40" />
                    <SPLIT distance="300" swimtime="00:03:28.82" />
                    <SPLIT distance="325" swimtime="00:03:44.72" />
                    <SPLIT distance="350" swimtime="00:03:59.90" />
                    <SPLIT distance="375" swimtime="00:04:14.95" />
                    <SPLIT distance="400" swimtime="00:04:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="3" lane="7" heat="3" heatid="30036" swimtime="00:04:31.19" reactiontime="+72" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.51" />
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                    <SPLIT distance="75" swimtime="00:00:46.36" />
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                    <SPLIT distance="125" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:01:37.53" />
                    <SPLIT distance="175" swimtime="00:01:54.60" />
                    <SPLIT distance="200" swimtime="00:02:11.31" />
                    <SPLIT distance="225" swimtime="00:02:30.72" />
                    <SPLIT distance="250" swimtime="00:02:50.18" />
                    <SPLIT distance="275" swimtime="00:03:09.79" />
                    <SPLIT distance="300" swimtime="00:03:29.64" />
                    <SPLIT distance="325" swimtime="00:03:45.70" />
                    <SPLIT distance="350" swimtime="00:04:01.18" />
                    <SPLIT distance="375" swimtime="00:04:16.36" />
                    <SPLIT distance="400" swimtime="00:04:31.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="171067" lastname="NAMBA" firstname="Miyu" gender="F" birthdate="2002-05-31">
              <ENTRIES>
                <ENTRY entrytime="00:03:59.47" eventid="1" heat="4" lane="5">
                  <MEETINFO date="2021-10-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:08:15.47" eventid="12" heat="0" lane="2147483647">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="00:16:12.97" eventid="33" heat="0" lane="-1">
                  <MEETINFO date="2022-03-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="101" place="4" lane="2" heat="1" heatid="10101" swimtime="00:04:01.13" reactiontime="+75" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="75" swimtime="00:00:43.22" />
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                    <SPLIT distance="125" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:28.91" />
                    <SPLIT distance="175" swimtime="00:01:44.15" />
                    <SPLIT distance="200" swimtime="00:01:59.50" />
                    <SPLIT distance="225" swimtime="00:02:14.81" />
                    <SPLIT distance="250" swimtime="00:02:30.27" />
                    <SPLIT distance="275" swimtime="00:02:45.70" />
                    <SPLIT distance="300" swimtime="00:03:01.11" />
                    <SPLIT distance="325" swimtime="00:03:16.26" />
                    <SPLIT distance="350" swimtime="00:03:31.36" />
                    <SPLIT distance="375" swimtime="00:03:46.49" />
                    <SPLIT distance="400" swimtime="00:04:01.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="5" lane="5" heat="4" heatid="40001" swimtime="00:04:00.97" reactiontime="+69" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:00:57.46" />
                    <SPLIT distance="125" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:27.45" />
                    <SPLIT distance="175" swimtime="00:01:42.58" />
                    <SPLIT distance="200" swimtime="00:01:58.05" />
                    <SPLIT distance="225" swimtime="00:02:13.54" />
                    <SPLIT distance="250" swimtime="00:02:29.08" />
                    <SPLIT distance="275" swimtime="00:02:44.56" />
                    <SPLIT distance="300" swimtime="00:03:00.12" />
                    <SPLIT distance="325" swimtime="00:03:15.38" />
                    <SPLIT distance="350" swimtime="00:03:30.90" />
                    <SPLIT distance="375" swimtime="00:03:46.25" />
                    <SPLIT distance="400" swimtime="00:04:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="3" lane="6" heat="5" heatid="30112" swimtime="00:08:12.98" reactiontime="+71" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="75" swimtime="00:00:44.12" />
                    <SPLIT distance="100" swimtime="00:00:59.59" />
                    <SPLIT distance="125" swimtime="00:01:14.98" />
                    <SPLIT distance="150" swimtime="00:01:30.51" />
                    <SPLIT distance="175" swimtime="00:01:45.95" />
                    <SPLIT distance="200" swimtime="00:02:01.38" />
                    <SPLIT distance="225" swimtime="00:02:16.84" />
                    <SPLIT distance="250" swimtime="00:02:32.45" />
                    <SPLIT distance="275" swimtime="00:02:48.02" />
                    <SPLIT distance="300" swimtime="00:03:03.72" />
                    <SPLIT distance="325" swimtime="00:03:19.33" />
                    <SPLIT distance="350" swimtime="00:03:34.94" />
                    <SPLIT distance="375" swimtime="00:03:50.45" />
                    <SPLIT distance="400" swimtime="00:04:06.20" />
                    <SPLIT distance="425" swimtime="00:04:21.81" />
                    <SPLIT distance="450" swimtime="00:04:37.53" />
                    <SPLIT distance="475" swimtime="00:04:53.18" />
                    <SPLIT distance="500" swimtime="00:05:08.70" />
                    <SPLIT distance="525" swimtime="00:05:24.48" />
                    <SPLIT distance="550" swimtime="00:05:40.15" />
                    <SPLIT distance="575" swimtime="00:05:55.66" />
                    <SPLIT distance="600" swimtime="00:06:11.33" />
                    <SPLIT distance="625" swimtime="00:06:26.82" />
                    <SPLIT distance="650" swimtime="00:06:42.40" />
                    <SPLIT distance="675" swimtime="00:06:57.86" />
                    <SPLIT distance="700" swimtime="00:07:13.54" />
                    <SPLIT distance="725" swimtime="00:07:28.80" />
                    <SPLIT distance="750" swimtime="00:07:44.14" />
                    <SPLIT distance="775" swimtime="00:07:58.80" />
                    <SPLIT distance="800" swimtime="00:08:12.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="2" lane="8" heat="5" heatid="30133" swimtime="00:15:46.76" reactiontime="+75" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                    <SPLIT distance="75" swimtime="00:00:44.99" />
                    <SPLIT distance="100" swimtime="00:01:00.80" />
                    <SPLIT distance="125" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:01:32.43" />
                    <SPLIT distance="175" swimtime="00:01:48.31" />
                    <SPLIT distance="200" swimtime="00:02:04.22" />
                    <SPLIT distance="225" swimtime="00:02:20.17" />
                    <SPLIT distance="250" swimtime="00:02:36.00" />
                    <SPLIT distance="275" swimtime="00:02:51.84" />
                    <SPLIT distance="300" swimtime="00:03:07.74" />
                    <SPLIT distance="325" swimtime="00:03:23.61" />
                    <SPLIT distance="350" swimtime="00:03:39.32" />
                    <SPLIT distance="375" swimtime="00:03:55.07" />
                    <SPLIT distance="400" swimtime="00:04:10.86" />
                    <SPLIT distance="425" swimtime="00:04:26.73" />
                    <SPLIT distance="450" swimtime="00:04:42.49" />
                    <SPLIT distance="475" swimtime="00:04:58.35" />
                    <SPLIT distance="500" swimtime="00:05:14.10" />
                    <SPLIT distance="525" swimtime="00:05:30.01" />
                    <SPLIT distance="550" swimtime="00:05:45.78" />
                    <SPLIT distance="575" swimtime="00:06:01.58" />
                    <SPLIT distance="600" swimtime="00:06:17.48" />
                    <SPLIT distance="625" swimtime="00:06:33.30" />
                    <SPLIT distance="650" swimtime="00:06:49.17" />
                    <SPLIT distance="675" swimtime="00:07:04.97" />
                    <SPLIT distance="700" swimtime="00:07:20.82" />
                    <SPLIT distance="725" swimtime="00:07:36.78" />
                    <SPLIT distance="750" swimtime="00:07:52.68" />
                    <SPLIT distance="775" swimtime="00:08:08.67" />
                    <SPLIT distance="800" swimtime="00:08:24.60" />
                    <SPLIT distance="825" swimtime="00:08:40.56" />
                    <SPLIT distance="850" swimtime="00:08:56.42" />
                    <SPLIT distance="875" swimtime="00:09:12.37" />
                    <SPLIT distance="900" swimtime="00:09:28.31" />
                    <SPLIT distance="925" swimtime="00:09:44.22" />
                    <SPLIT distance="950" swimtime="00:10:00.08" />
                    <SPLIT distance="975" swimtime="00:10:16.06" />
                    <SPLIT distance="1000" swimtime="00:10:32.02" />
                    <SPLIT distance="1025" swimtime="00:10:47.83" />
                    <SPLIT distance="1050" swimtime="00:11:03.80" />
                    <SPLIT distance="1075" swimtime="00:11:19.84" />
                    <SPLIT distance="1100" swimtime="00:11:35.75" />
                    <SPLIT distance="1125" swimtime="00:11:51.75" />
                    <SPLIT distance="1150" swimtime="00:12:07.76" />
                    <SPLIT distance="1175" swimtime="00:12:23.66" />
                    <SPLIT distance="1200" swimtime="00:12:39.70" />
                    <SPLIT distance="1225" swimtime="00:12:55.72" />
                    <SPLIT distance="1250" swimtime="00:13:11.65" />
                    <SPLIT distance="1275" swimtime="00:13:27.59" />
                    <SPLIT distance="1300" swimtime="00:13:43.56" />
                    <SPLIT distance="1325" swimtime="00:13:59.57" />
                    <SPLIT distance="1350" swimtime="00:14:15.52" />
                    <SPLIT distance="1375" swimtime="00:14:31.39" />
                    <SPLIT distance="1400" swimtime="00:14:47.10" />
                    <SPLIT distance="1425" swimtime="00:15:02.71" />
                    <SPLIT distance="1450" swimtime="00:15:18.06" />
                    <SPLIT distance="1475" swimtime="00:15:32.75" />
                    <SPLIT distance="1500" swimtime="00:15:46.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210166" lastname="SUZUKI" firstname="Ayami" gender="F" birthdate="2005-05-13">
              <ENTRIES>
                <ENTRY entrytime="00:04:32.02" eventid="36" heat="4" lane="2">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="36" place="16" lane="2" heat="4" heatid="40036" swimtime="00:04:40.95" reactiontime="+56" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="75" swimtime="00:00:44.70" />
                    <SPLIT distance="100" swimtime="00:01:01.35" />
                    <SPLIT distance="125" swimtime="00:01:18.73" />
                    <SPLIT distance="150" swimtime="00:01:35.52" />
                    <SPLIT distance="175" swimtime="00:01:52.67" />
                    <SPLIT distance="200" swimtime="00:02:09.85" />
                    <SPLIT distance="225" swimtime="00:02:30.51" />
                    <SPLIT distance="250" swimtime="00:02:51.12" />
                    <SPLIT distance="275" swimtime="00:03:12.19" />
                    <SPLIT distance="300" swimtime="00:03:33.29" />
                    <SPLIT distance="325" swimtime="00:03:50.62" />
                    <SPLIT distance="350" swimtime="00:04:07.57" />
                    <SPLIT distance="375" swimtime="00:04:24.44" />
                    <SPLIT distance="400" swimtime="00:04:40.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130475" lastname="TAKAHASHI" firstname="Miki" gender="F" birthdate="1995-04-10">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:26.55" eventid="18" heat="6" lane="7">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="19" lane="7" heat="6" heatid="60018" swimtime="00:00:26.77" reactiontime="+56" points="841">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214396" lastname="JINNO" firstname="Yume" gender="F" birthdate="2002-11-23">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:24.49" eventid="30" heat="7" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="30" place="18" lane="7" heat="7" heatid="70030" swimtime="00:00:24.74" reactiontime="+58" points="796">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:24.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141380" lastname="MORIYAMA" firstname="Yukimi" gender="F" birthdate="1996-08-09">
              <ENTRIES>
                <ENTRY entrytime="00:08:24.83" eventid="12" heat="2" lane="4">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="9" lane="4" heat="2" heatid="20012" swimtime="00:08:25.46" reactiontime="+68" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                    <SPLIT distance="75" swimtime="00:00:44.35" />
                    <SPLIT distance="100" swimtime="00:01:00.17" />
                    <SPLIT distance="125" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:31.89" />
                    <SPLIT distance="175" swimtime="00:01:47.86" />
                    <SPLIT distance="200" swimtime="00:02:03.85" />
                    <SPLIT distance="225" swimtime="00:02:19.80" />
                    <SPLIT distance="250" swimtime="00:02:35.68" />
                    <SPLIT distance="275" swimtime="00:02:51.67" />
                    <SPLIT distance="300" swimtime="00:03:07.37" />
                    <SPLIT distance="325" swimtime="00:03:23.70" />
                    <SPLIT distance="350" swimtime="00:03:39.66" />
                    <SPLIT distance="375" swimtime="00:03:55.85" />
                    <SPLIT distance="400" swimtime="00:04:11.80" />
                    <SPLIT distance="425" swimtime="00:04:27.82" />
                    <SPLIT distance="450" swimtime="00:04:43.92" />
                    <SPLIT distance="475" swimtime="00:05:00.08" />
                    <SPLIT distance="500" swimtime="00:05:16.09" />
                    <SPLIT distance="525" swimtime="00:05:32.17" />
                    <SPLIT distance="550" swimtime="00:05:48.17" />
                    <SPLIT distance="575" swimtime="00:06:04.09" />
                    <SPLIT distance="600" swimtime="00:06:19.88" />
                    <SPLIT distance="625" swimtime="00:06:36.11" />
                    <SPLIT distance="650" swimtime="00:06:52.26" />
                    <SPLIT distance="675" swimtime="00:07:08.21" />
                    <SPLIT distance="700" swimtime="00:07:24.22" />
                    <SPLIT distance="725" swimtime="00:07:40.14" />
                    <SPLIT distance="750" swimtime="00:07:56.04" />
                    <SPLIT distance="775" swimtime="00:08:11.41" />
                    <SPLIT distance="800" swimtime="00:08:25.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214524" lastname="MATSUMOTO" firstname="Shuya" gender="M" birthdate="2000-05-10">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:52.17" eventid="23" heat="3" lane="6">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="23" place="4" lane="6" heat="3" heatid="30023" swimtime="00:00:51.99" reactiontime="+61" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:23.28" />
                    <SPLIT distance="75" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="9" lane="5" heat="1" heatid="10223" swimtime="00:00:51.99" reactiontime="+59" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.52" />
                    <SPLIT distance="50" swimtime="00:00:23.05" />
                    <SPLIT distance="75" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214395" lastname="WATANABE" firstname="Temma" gender="M" birthdate="2002-09-11" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Japan">
              <RESULTS>
                <RESULT eventid="109" place="7" lane="8" heat="1" swimtime="00:03:07.93" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.47" />
                    <SPLIT distance="75" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:00:46.72" />
                    <SPLIT distance="125" swimtime="00:00:56.76" />
                    <SPLIT distance="150" swimtime="00:01:08.66" />
                    <SPLIT distance="175" swimtime="00:01:20.97" />
                    <SPLIT distance="200" swimtime="00:01:33.35" />
                    <SPLIT distance="225" swimtime="00:01:43.55" />
                    <SPLIT distance="250" swimtime="00:01:55.45" />
                    <SPLIT distance="275" swimtime="00:02:07.93" />
                    <SPLIT distance="300" swimtime="00:02:20.28" />
                    <SPLIT distance="325" swimtime="00:02:30.83" />
                    <SPLIT distance="350" swimtime="00:02:43.00" />
                    <SPLIT distance="375" swimtime="00:02:55.57" />
                    <SPLIT distance="400" swimtime="00:03:07.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130459" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="108761" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="214380" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="214381" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="8" lane="2" heat="2" swimtime="00:03:09.25" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.99" />
                    <SPLIT distance="50" swimtime="00:00:22.96" />
                    <SPLIT distance="75" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:00:47.90" />
                    <SPLIT distance="125" swimtime="00:00:58.16" />
                    <SPLIT distance="150" swimtime="00:01:10.17" />
                    <SPLIT distance="175" swimtime="00:01:22.52" />
                    <SPLIT distance="200" swimtime="00:01:34.67" />
                    <SPLIT distance="225" swimtime="00:01:44.79" />
                    <SPLIT distance="250" swimtime="00:01:56.71" />
                    <SPLIT distance="275" swimtime="00:02:09.16" />
                    <SPLIT distance="300" swimtime="00:02:21.62" />
                    <SPLIT distance="325" swimtime="00:02:32.16" />
                    <SPLIT distance="350" swimtime="00:02:44.30" />
                    <SPLIT distance="375" swimtime="00:02:56.88" />
                    <SPLIT distance="400" swimtime="00:03:09.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130459" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="108761" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="214380" reactiontime="+15" />
                    <RELAYPOSITION number="4" athleteid="214381" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Japan">
              <RESULTS>
                <RESULT eventid="148" place="4" lane="5" heat="1" swimtime="00:03:22.70" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                    <SPLIT distance="75" swimtime="00:00:36.83" />
                    <SPLIT distance="100" swimtime="00:00:49.98" />
                    <SPLIT distance="125" swimtime="00:01:01.67" />
                    <SPLIT distance="150" swimtime="00:01:15.97" />
                    <SPLIT distance="175" swimtime="00:01:30.79" />
                    <SPLIT distance="200" swimtime="00:01:46.25" />
                    <SPLIT distance="225" swimtime="00:01:56.82" />
                    <SPLIT distance="250" swimtime="00:02:09.40" />
                    <SPLIT distance="275" swimtime="00:02:22.42" />
                    <SPLIT distance="300" swimtime="00:02:36.31" />
                    <SPLIT distance="325" swimtime="00:02:46.60" />
                    <SPLIT distance="350" swimtime="00:02:58.50" />
                    <SPLIT distance="375" swimtime="00:03:10.68" />
                    <SPLIT distance="400" swimtime="00:03:22.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101144" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="191038" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="149684" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="130459" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="2" lane="6" heat="2" swimtime="00:03:23.68" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                    <SPLIT distance="75" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:00:50.43" />
                    <SPLIT distance="125" swimtime="00:01:02.06" />
                    <SPLIT distance="150" swimtime="00:01:16.60" />
                    <SPLIT distance="175" swimtime="00:01:31.51" />
                    <SPLIT distance="200" swimtime="00:01:46.92" />
                    <SPLIT distance="225" swimtime="00:01:57.28" />
                    <SPLIT distance="250" swimtime="00:02:10.03" />
                    <SPLIT distance="275" swimtime="00:02:23.23" />
                    <SPLIT distance="300" swimtime="00:02:36.98" />
                    <SPLIT distance="325" swimtime="00:02:47.16" />
                    <SPLIT distance="350" swimtime="00:02:59.05" />
                    <SPLIT distance="375" swimtime="00:03:11.37" />
                    <SPLIT distance="400" swimtime="00:03:23.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101144" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="129138" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="214386" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="108761" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Japan">
              <RESULTS>
                <RESULT eventid="132" place="5" lane="5" heat="1" swimtime="00:06:52.04" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.08" />
                    <SPLIT distance="50" swimtime="00:00:23.75" />
                    <SPLIT distance="75" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:00:49.85" />
                    <SPLIT distance="125" swimtime="00:01:03.35" />
                    <SPLIT distance="150" swimtime="00:01:16.84" />
                    <SPLIT distance="175" swimtime="00:01:30.57" />
                    <SPLIT distance="200" swimtime="00:01:43.78" />
                    <SPLIT distance="225" swimtime="00:01:54.05" />
                    <SPLIT distance="250" swimtime="00:02:06.16" />
                    <SPLIT distance="275" swimtime="00:02:18.79" />
                    <SPLIT distance="300" swimtime="00:02:31.71" />
                    <SPLIT distance="325" swimtime="00:02:44.91" />
                    <SPLIT distance="350" swimtime="00:02:58.15" />
                    <SPLIT distance="375" swimtime="00:03:11.42" />
                    <SPLIT distance="400" swimtime="00:03:24.44" />
                    <SPLIT distance="425" swimtime="00:03:35.17" />
                    <SPLIT distance="450" swimtime="00:03:47.68" />
                    <SPLIT distance="475" swimtime="00:04:00.40" />
                    <SPLIT distance="500" swimtime="00:04:13.35" />
                    <SPLIT distance="525" swimtime="00:04:26.77" />
                    <SPLIT distance="550" swimtime="00:04:40.25" />
                    <SPLIT distance="575" swimtime="00:04:54.15" />
                    <SPLIT distance="600" swimtime="00:05:07.62" />
                    <SPLIT distance="625" swimtime="00:05:18.15" />
                    <SPLIT distance="650" swimtime="00:05:30.71" />
                    <SPLIT distance="675" swimtime="00:05:43.68" />
                    <SPLIT distance="700" swimtime="00:05:57.17" />
                    <SPLIT distance="725" swimtime="00:06:10.73" />
                    <SPLIT distance="750" swimtime="00:06:24.64" />
                    <SPLIT distance="775" swimtime="00:06:38.51" />
                    <SPLIT distance="800" swimtime="00:06:52.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214395" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="130459" reactiontime="+9" />
                    <RELAYPOSITION number="3" athleteid="214381" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="214524" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="2" lane="6" heat="2" swimtime="00:06:54.26" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.14" />
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                    <SPLIT distance="75" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:00:49.85" />
                    <SPLIT distance="125" swimtime="00:01:03.11" />
                    <SPLIT distance="150" swimtime="00:01:16.63" />
                    <SPLIT distance="175" swimtime="00:01:30.25" />
                    <SPLIT distance="200" swimtime="00:01:43.45" />
                    <SPLIT distance="225" swimtime="00:01:54.47" />
                    <SPLIT distance="250" swimtime="00:02:07.17" />
                    <SPLIT distance="275" swimtime="00:02:20.23" />
                    <SPLIT distance="300" swimtime="00:02:33.41" />
                    <SPLIT distance="325" swimtime="00:02:46.68" />
                    <SPLIT distance="350" swimtime="00:03:00.27" />
                    <SPLIT distance="375" swimtime="00:03:13.93" />
                    <SPLIT distance="400" swimtime="00:03:27.04" />
                    <SPLIT distance="425" swimtime="00:03:38.08" />
                    <SPLIT distance="450" swimtime="00:03:51.04" />
                    <SPLIT distance="475" swimtime="00:04:04.20" />
                    <SPLIT distance="500" swimtime="00:04:17.44" />
                    <SPLIT distance="525" swimtime="00:04:30.68" />
                    <SPLIT distance="550" swimtime="00:04:44.14" />
                    <SPLIT distance="575" swimtime="00:04:57.96" />
                    <SPLIT distance="600" swimtime="00:05:11.63" />
                    <SPLIT distance="625" swimtime="00:05:22.31" />
                    <SPLIT distance="650" swimtime="00:05:34.85" />
                    <SPLIT distance="675" swimtime="00:05:47.69" />
                    <SPLIT distance="700" swimtime="00:06:01.04" />
                    <SPLIT distance="725" swimtime="00:06:14.39" />
                    <SPLIT distance="750" swimtime="00:06:27.81" />
                    <SPLIT distance="775" swimtime="00:06:41.20" />
                    <SPLIT distance="800" swimtime="00:06:54.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214395" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="214381" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="214524" reactiontime="+49" />
                    <RELAYPOSITION number="4" athleteid="130459" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Japan">
              <RESULTS>
                <RESULT eventid="126" place="4" lane="6" heat="1" swimtime="00:01:23.80" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.03" />
                    <SPLIT distance="50" swimtime="00:00:21.26" />
                    <SPLIT distance="75" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:00:42.05" />
                    <SPLIT distance="125" swimtime="00:00:51.71" />
                    <SPLIT distance="150" swimtime="00:01:02.84" />
                    <SPLIT distance="175" swimtime="00:01:12.65" />
                    <SPLIT distance="200" swimtime="00:01:23.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130485" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="214380" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="118529" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="108761" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="4" lane="2" heat="1" swimtime="00:01:24.17" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.02" />
                    <SPLIT distance="50" swimtime="00:00:21.14" />
                    <SPLIT distance="75" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:00:42.03" />
                    <SPLIT distance="125" swimtime="00:00:51.98" />
                    <SPLIT distance="150" swimtime="00:01:03.09" />
                    <SPLIT distance="175" swimtime="00:01:12.98" />
                    <SPLIT distance="200" swimtime="00:01:24.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130485" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="214380" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="118529" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="108761" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Japan">
              <RESULTS>
                <RESULT eventid="127" place="5" lane="1" heat="1" swimtime="00:01:30.05" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.98" />
                    <SPLIT distance="50" swimtime="00:00:21.24" />
                    <SPLIT distance="75" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:00:42.05" />
                    <SPLIT distance="125" swimtime="00:00:53.30" />
                    <SPLIT distance="150" swimtime="00:01:06.07" />
                    <SPLIT distance="175" swimtime="00:01:17.41" />
                    <SPLIT distance="200" swimtime="00:01:30.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130485" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="214380" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="100703" reactiontime="+10" />
                    <RELAYPOSITION number="4" athleteid="153983" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="7" lane="6" heat="1" swimtime="00:01:31.49" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:21.57" />
                    <SPLIT distance="75" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:00:42.85" />
                    <SPLIT distance="125" swimtime="00:00:54.25" />
                    <SPLIT distance="150" swimtime="00:01:06.95" />
                    <SPLIT distance="175" swimtime="00:01:18.66" />
                    <SPLIT distance="200" swimtime="00:01:31.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214380" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="118529" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="100703" reactiontime="+4" />
                    <RELAYPOSITION number="4" athleteid="130475" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Japan">
              <RESULTS>
                <RESULT eventid="108" place="8" lane="8" heat="1" swimtime="00:03:34.78" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                    <SPLIT distance="75" swimtime="00:00:40.27" />
                    <SPLIT distance="100" swimtime="00:00:53.95" />
                    <SPLIT distance="125" swimtime="00:01:05.72" />
                    <SPLIT distance="150" swimtime="00:01:19.21" />
                    <SPLIT distance="175" swimtime="00:01:33.25" />
                    <SPLIT distance="200" swimtime="00:01:47.04" />
                    <SPLIT distance="225" swimtime="00:01:59.00" />
                    <SPLIT distance="250" swimtime="00:02:12.67" />
                    <SPLIT distance="275" swimtime="00:02:26.45" />
                    <SPLIT distance="300" swimtime="00:02:40.30" />
                    <SPLIT distance="325" swimtime="00:02:52.30" />
                    <SPLIT distance="350" swimtime="00:03:06.27" />
                    <SPLIT distance="375" swimtime="00:03:20.55" />
                    <SPLIT distance="400" swimtime="00:03:34.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="153984" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="100703" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="214396" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="130475" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="8" lane="6" heat="1" swimtime="00:03:33.64" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:25.97" />
                    <SPLIT distance="75" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:00:53.69" />
                    <SPLIT distance="125" swimtime="00:01:05.38" />
                    <SPLIT distance="150" swimtime="00:01:18.82" />
                    <SPLIT distance="175" swimtime="00:01:32.75" />
                    <SPLIT distance="200" swimtime="00:01:46.32" />
                    <SPLIT distance="225" swimtime="00:01:58.16" />
                    <SPLIT distance="250" swimtime="00:02:11.87" />
                    <SPLIT distance="275" swimtime="00:02:25.90" />
                    <SPLIT distance="300" swimtime="00:02:39.81" />
                    <SPLIT distance="325" swimtime="00:02:51.65" />
                    <SPLIT distance="350" swimtime="00:03:05.35" />
                    <SPLIT distance="375" swimtime="00:03:19.55" />
                    <SPLIT distance="400" swimtime="00:03:33.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="153984" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="100703" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="214396" reactiontime="+30" />
                    <RELAYPOSITION number="4" athleteid="130475" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Japan">
              <RESULTS>
                <RESULT eventid="147" place="-1" lane="2" heat="1" status="DSQ" swimtime="00:03:52.37" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                    <SPLIT distance="75" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:00:58.07" />
                    <SPLIT distance="125" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:28.20" />
                    <SPLIT distance="175" swimtime="00:01:45.09" />
                    <SPLIT distance="200" swimtime="00:02:02.72" />
                    <SPLIT distance="225" swimtime="00:02:14.65" />
                    <SPLIT distance="250" swimtime="00:02:29.00" />
                    <SPLIT distance="275" swimtime="00:02:44.13" />
                    <SPLIT distance="300" swimtime="00:02:59.91" />
                    <SPLIT distance="325" swimtime="00:03:11.21" />
                    <SPLIT distance="350" swimtime="00:03:24.69" />
                    <SPLIT distance="375" swimtime="00:03:38.60" />
                    <SPLIT distance="400" swimtime="00:03:52.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101276" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="130477" reactiontime="+38" />
                    <RELAYPOSITION number="3" athleteid="153983" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="100703" reactiontime="-7" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="5" lane="2" heat="2" swimtime="00:03:52.92" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="75" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:00:58.11" />
                    <SPLIT distance="125" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:28.05" />
                    <SPLIT distance="175" swimtime="00:01:45.03" />
                    <SPLIT distance="200" swimtime="00:02:02.42" />
                    <SPLIT distance="225" swimtime="00:02:14.45" />
                    <SPLIT distance="250" swimtime="00:02:29.02" />
                    <SPLIT distance="275" swimtime="00:02:43.97" />
                    <SPLIT distance="300" swimtime="00:02:59.40" />
                    <SPLIT distance="325" swimtime="00:03:11.31" />
                    <SPLIT distance="350" swimtime="00:03:24.85" />
                    <SPLIT distance="375" swimtime="00:03:38.92" />
                    <SPLIT distance="400" swimtime="00:03:52.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="153984" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="130477" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="153983" reactiontime="+45" />
                    <RELAYPOSITION number="4" athleteid="214396" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Japan">
              <RESULTS>
                <RESULT eventid="117" place="5" lane="1" heat="1" swimtime="00:07:44.87" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="75" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:00:56.20" />
                    <SPLIT distance="125" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:26.60" />
                    <SPLIT distance="175" swimtime="00:01:41.87" />
                    <SPLIT distance="200" swimtime="00:01:56.41" />
                    <SPLIT distance="225" swimtime="00:02:08.79" />
                    <SPLIT distance="250" swimtime="00:02:22.83" />
                    <SPLIT distance="275" swimtime="00:02:37.20" />
                    <SPLIT distance="300" swimtime="00:02:51.88" />
                    <SPLIT distance="325" swimtime="00:03:06.73" />
                    <SPLIT distance="350" swimtime="00:03:21.72" />
                    <SPLIT distance="375" swimtime="00:03:36.71" />
                    <SPLIT distance="400" swimtime="00:03:51.11" />
                    <SPLIT distance="425" swimtime="00:04:03.86" />
                    <SPLIT distance="450" swimtime="00:04:18.42" />
                    <SPLIT distance="475" swimtime="00:04:33.16" />
                    <SPLIT distance="500" swimtime="00:04:48.13" />
                    <SPLIT distance="525" swimtime="00:05:03.06" />
                    <SPLIT distance="550" swimtime="00:05:18.01" />
                    <SPLIT distance="575" swimtime="00:05:33.07" />
                    <SPLIT distance="600" swimtime="00:05:47.57" />
                    <SPLIT distance="625" swimtime="00:05:59.72" />
                    <SPLIT distance="650" swimtime="00:06:13.55" />
                    <SPLIT distance="675" swimtime="00:06:27.93" />
                    <SPLIT distance="700" swimtime="00:06:42.81" />
                    <SPLIT distance="725" swimtime="00:06:58.12" />
                    <SPLIT distance="750" swimtime="00:07:13.86" />
                    <SPLIT distance="775" swimtime="00:07:29.63" />
                    <SPLIT distance="800" swimtime="00:07:44.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100703" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="171067" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="149685" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="153984" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="7" lane="6" heat="1" swimtime="00:07:49.76" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.78" />
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                    <SPLIT distance="75" swimtime="00:00:42.16" />
                    <SPLIT distance="100" swimtime="00:00:57.26" />
                    <SPLIT distance="125" swimtime="00:01:12.47" />
                    <SPLIT distance="150" swimtime="00:01:27.75" />
                    <SPLIT distance="175" swimtime="00:01:42.80" />
                    <SPLIT distance="200" swimtime="00:01:57.05" />
                    <SPLIT distance="225" swimtime="00:02:09.86" />
                    <SPLIT distance="250" swimtime="00:02:24.59" />
                    <SPLIT distance="275" swimtime="00:02:39.40" />
                    <SPLIT distance="300" swimtime="00:02:54.35" />
                    <SPLIT distance="325" swimtime="00:03:09.35" />
                    <SPLIT distance="350" swimtime="00:03:24.39" />
                    <SPLIT distance="375" swimtime="00:03:39.41" />
                    <SPLIT distance="400" swimtime="00:03:53.86" />
                    <SPLIT distance="425" swimtime="00:04:06.67" />
                    <SPLIT distance="450" swimtime="00:04:21.25" />
                    <SPLIT distance="475" swimtime="00:04:35.95" />
                    <SPLIT distance="500" swimtime="00:04:51.03" />
                    <SPLIT distance="525" swimtime="00:05:05.79" />
                    <SPLIT distance="550" swimtime="00:05:20.94" />
                    <SPLIT distance="575" swimtime="00:05:35.80" />
                    <SPLIT distance="600" swimtime="00:05:50.55" />
                    <SPLIT distance="625" swimtime="00:06:03.43" />
                    <SPLIT distance="650" swimtime="00:06:18.22" />
                    <SPLIT distance="675" swimtime="00:06:33.11" />
                    <SPLIT distance="700" swimtime="00:06:48.28" />
                    <SPLIT distance="725" swimtime="00:07:03.64" />
                    <SPLIT distance="750" swimtime="00:07:19.21" />
                    <SPLIT distance="775" swimtime="00:07:34.76" />
                    <SPLIT distance="800" swimtime="00:07:49.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100703" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="171067" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="149685" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="153984" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Japan">
              <RESULTS>
                <RESULT eventid="125" place="7" lane="7" heat="1" swimtime="00:01:37.42" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:24.54" />
                    <SPLIT distance="75" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:00:48.97" />
                    <SPLIT distance="125" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:13.44" />
                    <SPLIT distance="175" swimtime="00:01:24.84" />
                    <SPLIT distance="200" swimtime="00:01:37.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100703" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="130475" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="214396" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="153983" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="6" lane="6" heat="2" swimtime="00:01:37.74" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:24.76" />
                    <SPLIT distance="75" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:00:49.09" />
                    <SPLIT distance="125" swimtime="00:01:00.65" />
                    <SPLIT distance="150" swimtime="00:01:13.44" />
                    <SPLIT distance="175" swimtime="00:01:24.89" />
                    <SPLIT distance="200" swimtime="00:01:37.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214396" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="130475" reactiontime="+4" />
                    <RELAYPOSITION number="3" athleteid="100703" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="153983" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Japan">
              <RESULTS>
                <RESULT eventid="134" place="7" lane="6" heat="1" swimtime="00:01:45.29" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                    <SPLIT distance="75" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:00:56.51" />
                    <SPLIT distance="125" swimtime="00:01:07.93" />
                    <SPLIT distance="150" swimtime="00:01:21.25" />
                    <SPLIT distance="175" swimtime="00:01:32.57" />
                    <SPLIT distance="200" swimtime="00:01:45.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130475" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="130477" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="214391" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="100703" reactiontime="+8" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="4" lane="1" heat="1" swimtime="00:01:45.41" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="75" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:00:56.24" />
                    <SPLIT distance="125" swimtime="00:01:07.44" />
                    <SPLIT distance="150" swimtime="00:01:20.97" />
                    <SPLIT distance="175" swimtime="00:01:32.58" />
                    <SPLIT distance="200" swimtime="00:01:45.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130475" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="130477" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="214391" reactiontime="+8" />
                    <RELAYPOSITION number="4" athleteid="214396" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Japan">
              <RESULTS>
                <RESULT eventid="111" place="6" lane="2" heat="1" swimtime="00:01:38.38" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                    <SPLIT distance="75" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:00:52.50" />
                    <SPLIT distance="125" swimtime="00:01:03.62" />
                    <SPLIT distance="150" swimtime="00:01:17.30" />
                    <SPLIT distance="175" swimtime="00:01:27.28" />
                    <SPLIT distance="200" swimtime="00:01:38.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130475" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="157430" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="153983" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="130485" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="5" lane="8" heat="4" swimtime="00:01:38.64" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                    <SPLIT distance="75" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:00:52.85" />
                    <SPLIT distance="125" swimtime="00:01:04.11" />
                    <SPLIT distance="150" swimtime="00:01:17.81" />
                    <SPLIT distance="175" swimtime="00:01:27.59" />
                    <SPLIT distance="200" swimtime="00:01:38.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130475" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="157430" reactiontime="+30" />
                    <RELAYPOSITION number="3" athleteid="214391" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="130485" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Japan">
              <RESULTS>
                <RESULT eventid="135" place="4" lane="6" heat="1" swimtime="00:01:31.28" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.18" />
                    <SPLIT distance="50" swimtime="00:00:22.93" />
                    <SPLIT distance="75" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:00:48.57" />
                    <SPLIT distance="125" swimtime="00:00:58.47" />
                    <SPLIT distance="150" swimtime="00:01:10.70" />
                    <SPLIT distance="175" swimtime="00:01:20.35" />
                    <SPLIT distance="200" swimtime="00:01:31.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="118529" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="191038" reactiontime="+3" />
                    <RELAYPOSITION number="3" athleteid="214386" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="214380" reactiontime="+10" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="4" lane="5" heat="2" swimtime="00:01:32.65" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:23.47" />
                    <SPLIT distance="75" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:00:49.41" />
                    <SPLIT distance="125" swimtime="00:00:59.53" />
                    <SPLIT distance="150" swimtime="00:01:11.60" />
                    <SPLIT distance="175" swimtime="00:01:21.46" />
                    <SPLIT distance="200" swimtime="00:01:32.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101144" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="191038" reactiontime="+14" />
                    <RELAYPOSITION number="3" athleteid="118529" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="130485" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Kazakhstan" shortname="KAZ" code="KAZ" nation="KAZ" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="137896" lastname="MUSSIN" firstname="Adilbek" gender="M" birthdate="1999-10-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.23" eventid="39" heat="5" lane="3">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.40" eventid="21" heat="2" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.50" eventid="5" heat="6" lane="7">
                  <MEETINFO date="2022-08-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="16" lane="3" heat="5" heatid="50039" swimtime="00:00:50.64" reactiontime="+69" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.88" />
                    <SPLIT distance="50" swimtime="00:00:23.83" />
                    <SPLIT distance="75" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:00:50.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="15" lane="8" heat="1" heatid="10239" swimtime="00:00:50.76" reactiontime="+68" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.85" />
                    <SPLIT distance="50" swimtime="00:00:23.63" />
                    <SPLIT distance="75" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:00:50.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="18" lane="7" heat="2" heatid="20021" swimtime="00:01:55.61" reactiontime="+69" points="820">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                    <SPLIT distance="75" swimtime="00:00:39.65" />
                    <SPLIT distance="100" swimtime="00:00:54.18" />
                    <SPLIT distance="125" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:23.91" />
                    <SPLIT distance="175" swimtime="00:01:39.34" />
                    <SPLIT distance="200" swimtime="00:01:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="32" lane="7" heat="6" heatid="60005" swimtime="00:00:23.09" reactiontime="+68" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.59" />
                    <SPLIT distance="50" swimtime="00:00:23.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153926" lastname="PCHELINTSEVA" firstname="Adelaida" gender="F" birthdate="1999-09-29">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.89" eventid="15" heat="3" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.62" eventid="40" heat="6" lane="8">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="37" lane="3" heat="3" heatid="30015" swimtime="00:01:09.42" reactiontime="+65" points="724">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="75" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:01:09.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="25" lane="8" heat="6" heatid="60040" swimtime="00:00:30.87" reactiontime="+63" points="791">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Kyrgyzstan" shortname="KGZ" code="KGZ" nation="KGZ" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="105376" lastname="PETRASHOV" firstname="Denis" gender="M" birthdate="2000-02-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.56" eventid="16" heat="5" lane="2">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.39" eventid="29" heat="4" lane="2">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.88" eventid="41" heat="7" lane="8">
                  <MEETINFO date="2021-10-08" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="24" lane="2" heat="5" heatid="50016" swimtime="00:00:58.21" reactiontime="+75" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="75" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:00:58.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="15" lane="2" heat="4" heatid="40029" swimtime="00:02:06.62" reactiontime="+79" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="75" swimtime="00:00:44.68" />
                    <SPLIT distance="100" swimtime="00:01:00.78" />
                    <SPLIT distance="125" swimtime="00:01:17.08" />
                    <SPLIT distance="150" swimtime="00:01:33.56" />
                    <SPLIT distance="175" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="21" lane="8" heat="7" heatid="70041" swimtime="00:00:26.71" reactiontime="+70" points="815">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Republic of Korea" shortname="KOR" code="KOR" nation="KOR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="145225" lastname="YANG" firstname="Jaehoon" gender="M" birthdate="1998-05-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.32" eventid="39" heat="4" lane="2">
                  <MEETINFO date="2022-03-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:00:22.85" eventid="31" heat="5" lane="5">
                  <MEETINFO date="2022-03-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="24" lane="2" heat="4" heatid="40039" swimtime="00:00:51.36" reactiontime="+67" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.83" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                    <SPLIT distance="75" swimtime="00:00:37.45" />
                    <SPLIT distance="100" swimtime="00:00:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="32" lane="5" heat="5" heatid="50031" swimtime="00:00:21.54" reactiontime="+67" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.37" />
                    <SPLIT distance="50" swimtime="00:00:21.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166111" lastname="HWANG" firstname="Sunwoo" gender="M" birthdate="2003-05-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.34" eventid="14" heat="9" lane="5">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.17" eventid="44" heat="4" lane="4">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="6" lane="5" heat="9" heatid="90014" swimtime="00:00:46.36" reactiontime="+63" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:22.18" />
                    <SPLIT distance="75" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="9" lane="3" heat="1" heatid="10214" swimtime="00:00:46.41" reactiontime="+61" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:22.44" />
                    <SPLIT distance="75" swimtime="00:00:34.51" />
                    <SPLIT distance="100" swimtime="00:00:46.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="144" place="1" lane="8" heat="1" heatid="10144" swimtime="00:01:39.72" reactiontime="+65" points="989">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.83" />
                    <SPLIT distance="50" swimtime="00:00:23.26" />
                    <SPLIT distance="75" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:00:48.88" />
                    <SPLIT distance="125" swimtime="00:01:01.46" />
                    <SPLIT distance="150" swimtime="00:01:14.20" />
                    <SPLIT distance="175" swimtime="00:01:27.00" />
                    <SPLIT distance="200" swimtime="00:01:39.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="8" lane="4" heat="4" heatid="40044" swimtime="00:01:42.44" reactiontime="+64" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:24.17" />
                    <SPLIT distance="75" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:00:50.51" />
                    <SPLIT distance="125" swimtime="00:01:03.56" />
                    <SPLIT distance="150" swimtime="00:01:16.74" />
                    <SPLIT distance="175" swimtime="00:01:30.00" />
                    <SPLIT distance="200" swimtime="00:01:42.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165487" lastname="KIM" firstname="Woomin" gender="M" birthdate="2001-08-24">
              <ENTRIES>
                <ENTRY entrytime="00:14:44.58" eventid="10" heat="2" lane="4">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:03:45.64" eventid="24" heat="3" lane="6">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:07:50.35" eventid="42" heat="2" lane="8">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="9" lane="4" heat="2" heatid="20010" swimtime="00:14:45.35" reactiontime="+59" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                    <SPLIT distance="75" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:00:54.07" />
                    <SPLIT distance="125" swimtime="00:01:08.07" />
                    <SPLIT distance="150" swimtime="00:01:22.32" />
                    <SPLIT distance="175" swimtime="00:01:36.66" />
                    <SPLIT distance="200" swimtime="00:01:50.92" />
                    <SPLIT distance="225" swimtime="00:02:05.28" />
                    <SPLIT distance="250" swimtime="00:02:19.74" />
                    <SPLIT distance="275" swimtime="00:02:34.09" />
                    <SPLIT distance="300" swimtime="00:02:48.57" />
                    <SPLIT distance="325" swimtime="00:03:03.02" />
                    <SPLIT distance="350" swimtime="00:03:17.44" />
                    <SPLIT distance="375" swimtime="00:03:31.91" />
                    <SPLIT distance="400" swimtime="00:03:46.32" />
                    <SPLIT distance="425" swimtime="00:04:00.66" />
                    <SPLIT distance="450" swimtime="00:04:15.17" />
                    <SPLIT distance="475" swimtime="00:04:29.73" />
                    <SPLIT distance="500" swimtime="00:04:44.36" />
                    <SPLIT distance="525" swimtime="00:04:59.05" />
                    <SPLIT distance="550" swimtime="00:05:13.69" />
                    <SPLIT distance="575" swimtime="00:05:28.32" />
                    <SPLIT distance="600" swimtime="00:05:42.96" />
                    <SPLIT distance="625" swimtime="00:05:57.65" />
                    <SPLIT distance="650" swimtime="00:06:12.38" />
                    <SPLIT distance="675" swimtime="00:06:27.23" />
                    <SPLIT distance="700" swimtime="00:06:42.02" />
                    <SPLIT distance="725" swimtime="00:06:56.87" />
                    <SPLIT distance="750" swimtime="00:07:11.73" />
                    <SPLIT distance="775" swimtime="00:07:26.56" />
                    <SPLIT distance="800" swimtime="00:07:41.42" />
                    <SPLIT distance="825" swimtime="00:07:56.27" />
                    <SPLIT distance="850" swimtime="00:08:11.22" />
                    <SPLIT distance="875" swimtime="00:08:26.09" />
                    <SPLIT distance="900" swimtime="00:08:41.18" />
                    <SPLIT distance="925" swimtime="00:08:56.28" />
                    <SPLIT distance="950" swimtime="00:09:11.38" />
                    <SPLIT distance="975" swimtime="00:09:26.55" />
                    <SPLIT distance="1000" swimtime="00:09:41.67" />
                    <SPLIT distance="1025" swimtime="00:09:56.87" />
                    <SPLIT distance="1050" swimtime="00:10:12.01" />
                    <SPLIT distance="1075" swimtime="00:10:27.27" />
                    <SPLIT distance="1100" swimtime="00:10:42.54" />
                    <SPLIT distance="1125" swimtime="00:10:57.95" />
                    <SPLIT distance="1150" swimtime="00:11:13.15" />
                    <SPLIT distance="1175" swimtime="00:11:28.30" />
                    <SPLIT distance="1200" swimtime="00:11:43.59" />
                    <SPLIT distance="1225" swimtime="00:11:59.01" />
                    <SPLIT distance="1250" swimtime="00:12:14.25" />
                    <SPLIT distance="1275" swimtime="00:12:29.61" />
                    <SPLIT distance="1300" swimtime="00:12:44.89" />
                    <SPLIT distance="1325" swimtime="00:13:00.03" />
                    <SPLIT distance="1350" swimtime="00:13:15.27" />
                    <SPLIT distance="1375" swimtime="00:13:30.43" />
                    <SPLIT distance="1400" swimtime="00:13:45.85" />
                    <SPLIT distance="1425" swimtime="00:14:01.01" />
                    <SPLIT distance="1450" swimtime="00:14:16.24" />
                    <SPLIT distance="1475" swimtime="00:14:31.32" />
                    <SPLIT distance="1500" swimtime="00:14:45.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="9" lane="6" heat="3" heatid="30024" swimtime="00:03:38.86" reactiontime="+58" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:24.52" />
                    <SPLIT distance="75" swimtime="00:00:38.11" />
                    <SPLIT distance="100" swimtime="00:00:51.79" />
                    <SPLIT distance="125" swimtime="00:01:05.52" />
                    <SPLIT distance="150" swimtime="00:01:19.42" />
                    <SPLIT distance="175" swimtime="00:01:33.38" />
                    <SPLIT distance="200" swimtime="00:01:47.39" />
                    <SPLIT distance="225" swimtime="00:02:01.23" />
                    <SPLIT distance="250" swimtime="00:02:15.28" />
                    <SPLIT distance="275" swimtime="00:02:29.32" />
                    <SPLIT distance="300" swimtime="00:02:43.43" />
                    <SPLIT distance="325" swimtime="00:02:57.53" />
                    <SPLIT distance="350" swimtime="00:03:11.53" />
                    <SPLIT distance="375" swimtime="00:03:25.39" />
                    <SPLIT distance="400" swimtime="00:03:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="12" lane="8" heat="2" heatid="20042" swimtime="00:07:45.29" reactiontime="+59" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="75" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:00:54.62" />
                    <SPLIT distance="125" swimtime="00:01:08.90" />
                    <SPLIT distance="150" swimtime="00:01:23.36" />
                    <SPLIT distance="175" swimtime="00:01:37.73" />
                    <SPLIT distance="200" swimtime="00:01:52.23" />
                    <SPLIT distance="225" swimtime="00:02:06.51" />
                    <SPLIT distance="250" swimtime="00:02:21.17" />
                    <SPLIT distance="275" swimtime="00:02:35.64" />
                    <SPLIT distance="300" swimtime="00:02:50.19" />
                    <SPLIT distance="325" swimtime="00:03:04.64" />
                    <SPLIT distance="350" swimtime="00:03:19.08" />
                    <SPLIT distance="375" swimtime="00:03:33.61" />
                    <SPLIT distance="400" swimtime="00:03:48.21" />
                    <SPLIT distance="425" swimtime="00:04:02.84" />
                    <SPLIT distance="450" swimtime="00:04:17.58" />
                    <SPLIT distance="475" swimtime="00:04:32.33" />
                    <SPLIT distance="500" swimtime="00:04:47.36" />
                    <SPLIT distance="525" swimtime="00:05:02.16" />
                    <SPLIT distance="550" swimtime="00:05:17.12" />
                    <SPLIT distance="575" swimtime="00:05:31.99" />
                    <SPLIT distance="600" swimtime="00:05:47.05" />
                    <SPLIT distance="625" swimtime="00:06:02.03" />
                    <SPLIT distance="650" swimtime="00:06:17.25" />
                    <SPLIT distance="675" swimtime="00:06:32.30" />
                    <SPLIT distance="700" swimtime="00:06:47.39" />
                    <SPLIT distance="725" swimtime="00:07:02.34" />
                    <SPLIT distance="750" swimtime="00:07:17.51" />
                    <SPLIT distance="775" swimtime="00:07:31.76" />
                    <SPLIT distance="800" swimtime="00:07:45.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214595" lastname="KIM" firstname="Sanha" gender="F" birthdate="1996-11-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.30" eventid="2" heat="3" lane="8">
                  <MEETINFO date="2022-03-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:28.68" eventid="18" heat="4" lane="2">
                  <MEETINFO date="2022-03-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="21" lane="8" heat="3" heatid="30002" swimtime="00:00:58.02" reactiontime="+53" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                    <SPLIT distance="75" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:00:58.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="18" lane="2" heat="4" heatid="40018" swimtime="00:00:26.70" reactiontime="+55" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:26.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201643" lastname="MOON" firstname="Sua" gender="F" birthdate="2008-11-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:08.50" eventid="15" heat="3" lane="5">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:26.64" eventid="28" heat="2" lane="2">
                  <MEETINFO date="2022-06-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="31" lane="5" heat="3" heatid="30015" swimtime="00:01:06.96" reactiontime="+64" points="807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="75" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="18" lane="2" heat="2" heatid="20028" swimtime="00:02:23.41" reactiontime="+63" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.17" />
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="75" swimtime="00:00:51.64" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="125" swimtime="00:01:28.58" />
                    <SPLIT distance="150" swimtime="00:01:46.83" />
                    <SPLIT distance="175" swimtime="00:02:05.20" />
                    <SPLIT distance="200" swimtime="00:02:23.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145245" lastname="KIM" firstname="Seoyeong" gender="F" birthdate="1994-03-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.32" eventid="38" heat="2" lane="1">
                  <MEETINFO date="2022-03-24" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.60" eventid="6" heat="4" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="13" lane="1" heat="2" heatid="20038" swimtime="00:00:57.26" reactiontime="+56" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="75" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:00:57.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="11" lane="1" heat="2" heatid="20238" swimtime="00:00:57.07" reactiontime="+54" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.26" />
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                    <SPLIT distance="75" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:00:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="11" lane="2" heat="4" heatid="40006" swimtime="00:02:07.74" reactiontime="+62" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                    <SPLIT distance="75" swimtime="00:00:43.55" />
                    <SPLIT distance="100" swimtime="00:00:59.02" />
                    <SPLIT distance="125" swimtime="00:01:17.62" />
                    <SPLIT distance="150" swimtime="00:01:36.64" />
                    <SPLIT distance="175" swimtime="00:01:52.60" />
                    <SPLIT distance="200" swimtime="00:02:07.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201667" lastname="HUR" firstname="Yeonkyung" gender="F" birthdate="2005-12-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.22" eventid="13" heat="6" lane="8">
                  <MEETINFO date="2022-03-25" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.27" eventid="43" heat="2" lane="2">
                  <MEETINFO date="2022-03-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:25.70" eventid="30" heat="5" lane="1">
                  <MEETINFO date="2022-03-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="32" lane="8" heat="6" heatid="60013" swimtime="00:00:54.59" reactiontime="+70" points="779">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                    <SPLIT distance="75" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:00:54.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="21" lane="2" heat="2" heatid="20043" swimtime="00:01:58.41" reactiontime="+66" points="808">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                    <SPLIT distance="75" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="125" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:29.01" />
                    <SPLIT distance="175" swimtime="00:01:44.23" />
                    <SPLIT distance="200" swimtime="00:01:58.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="24" lane="1" heat="5" heatid="50030" swimtime="00:00:24.99" reactiontime="+66" points="772">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154128" lastname="LEE" firstname="Hojoon" gender="M" birthdate="2001-02-14" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Republic of Korea">
              <RESULTS>
                <RESULT eventid="132" place="4" lane="2" heat="1" swimtime="00:06:49.67" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.85" />
                    <SPLIT distance="50" swimtime="00:00:23.33" />
                    <SPLIT distance="75" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:00:48.79" />
                    <SPLIT distance="125" swimtime="00:01:01.77" />
                    <SPLIT distance="150" swimtime="00:01:14.97" />
                    <SPLIT distance="175" swimtime="00:01:28.24" />
                    <SPLIT distance="200" swimtime="00:01:40.99" />
                    <SPLIT distance="225" swimtime="00:01:51.57" />
                    <SPLIT distance="250" swimtime="00:02:04.06" />
                    <SPLIT distance="275" swimtime="00:02:16.82" />
                    <SPLIT distance="300" swimtime="00:02:29.83" />
                    <SPLIT distance="325" swimtime="00:02:42.93" />
                    <SPLIT distance="350" swimtime="00:02:56.27" />
                    <SPLIT distance="375" swimtime="00:03:09.69" />
                    <SPLIT distance="400" swimtime="00:03:23.02" />
                    <SPLIT distance="425" swimtime="00:03:34.13" />
                    <SPLIT distance="450" swimtime="00:03:46.95" />
                    <SPLIT distance="475" swimtime="00:03:59.86" />
                    <SPLIT distance="500" swimtime="00:04:12.88" />
                    <SPLIT distance="525" swimtime="00:04:25.98" />
                    <SPLIT distance="550" swimtime="00:04:39.33" />
                    <SPLIT distance="575" swimtime="00:04:52.81" />
                    <SPLIT distance="600" swimtime="00:05:05.94" />
                    <SPLIT distance="625" swimtime="00:05:16.46" />
                    <SPLIT distance="650" swimtime="00:05:29.16" />
                    <SPLIT distance="675" swimtime="00:05:42.09" />
                    <SPLIT distance="700" swimtime="00:05:55.30" />
                    <SPLIT distance="725" swimtime="00:06:08.73" />
                    <SPLIT distance="750" swimtime="00:06:22.47" />
                    <SPLIT distance="775" swimtime="00:06:36.37" />
                    <SPLIT distance="800" swimtime="00:06:49.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="166111" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="165487" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="154128" reactiontime="+33" />
                    <RELAYPOSITION number="4" athleteid="145225" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="5" lane="3" heat="1" swimtime="00:06:55.24" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.11" />
                    <SPLIT distance="50" swimtime="00:00:23.68" />
                    <SPLIT distance="75" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:00:49.47" />
                    <SPLIT distance="125" swimtime="00:01:02.39" />
                    <SPLIT distance="150" swimtime="00:01:15.52" />
                    <SPLIT distance="175" swimtime="00:01:28.87" />
                    <SPLIT distance="200" swimtime="00:01:41.97" />
                    <SPLIT distance="225" swimtime="00:01:52.76" />
                    <SPLIT distance="250" swimtime="00:02:05.32" />
                    <SPLIT distance="275" swimtime="00:02:18.14" />
                    <SPLIT distance="300" swimtime="00:02:31.32" />
                    <SPLIT distance="325" swimtime="00:02:44.72" />
                    <SPLIT distance="350" swimtime="00:02:58.17" />
                    <SPLIT distance="375" swimtime="00:03:11.76" />
                    <SPLIT distance="400" swimtime="00:03:24.92" />
                    <SPLIT distance="425" swimtime="00:03:36.05" />
                    <SPLIT distance="450" swimtime="00:03:48.71" />
                    <SPLIT distance="475" swimtime="00:04:01.79" />
                    <SPLIT distance="500" swimtime="00:04:15.04" />
                    <SPLIT distance="525" swimtime="00:04:28.33" />
                    <SPLIT distance="550" swimtime="00:04:41.80" />
                    <SPLIT distance="575" swimtime="00:04:55.41" />
                    <SPLIT distance="600" swimtime="00:05:08.49" />
                    <SPLIT distance="625" swimtime="00:05:19.70" />
                    <SPLIT distance="650" swimtime="00:05:32.74" />
                    <SPLIT distance="675" swimtime="00:05:46.17" />
                    <SPLIT distance="700" swimtime="00:05:59.66" />
                    <SPLIT distance="725" swimtime="00:06:13.41" />
                    <SPLIT distance="750" swimtime="00:06:27.19" />
                    <SPLIT distance="775" swimtime="00:06:41.43" />
                    <SPLIT distance="800" swimtime="00:06:55.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="166111" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="165487" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="154128" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="145225" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Republic of Korea">
              <RESULTS>
                <RESULT eventid="47" place="10" lane="7" heat="1" swimtime="00:03:56.66" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:27.64" />
                    <SPLIT distance="75" swimtime="00:00:42.80" />
                    <SPLIT distance="100" swimtime="00:00:58.01" />
                    <SPLIT distance="125" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:29.24" />
                    <SPLIT distance="175" swimtime="00:01:46.87" />
                    <SPLIT distance="200" swimtime="00:02:04.88" />
                    <SPLIT distance="225" swimtime="00:02:16.88" />
                    <SPLIT distance="250" swimtime="00:02:31.48" />
                    <SPLIT distance="275" swimtime="00:02:46.69" />
                    <SPLIT distance="300" swimtime="00:03:02.67" />
                    <SPLIT distance="325" swimtime="00:03:14.75" />
                    <SPLIT distance="350" swimtime="00:03:28.63" />
                    <SPLIT distance="375" swimtime="00:03:42.96" />
                    <SPLIT distance="400" swimtime="00:03:56.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214595" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="201643" reactiontime="+5" />
                    <RELAYPOSITION number="3" athleteid="145245" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="201667" reactiontime="+6" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Republic of Korea">
              <RESULTS>
                <RESULT eventid="34" place="9" lane="1" heat="2" swimtime="00:01:48.24" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.03" />
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                    <SPLIT distance="75" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:00:57.85" />
                    <SPLIT distance="125" swimtime="00:01:09.41" />
                    <SPLIT distance="150" swimtime="00:01:23.68" />
                    <SPLIT distance="175" swimtime="00:01:35.53" />
                    <SPLIT distance="200" swimtime="00:01:48.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214595" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="201643" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="145245" reactiontime="+3" />
                    <RELAYPOSITION number="4" athleteid="201667" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Kosovo" shortname="KOS" code="KOS" nation="KOS" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="198067" lastname="MUJA" firstname="Martin" gender="M" birthdate="2004-07-22">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.30" eventid="14" heat="3" lane="8">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.61" eventid="31" heat="4" lane="6">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="65" lane="8" heat="3" heatid="30014" swimtime="00:00:52.28" reactiontime="+65" points="630">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.57" />
                    <SPLIT distance="50" swimtime="00:00:24.59" />
                    <SPLIT distance="75" swimtime="00:00:38.17" />
                    <SPLIT distance="100" swimtime="00:00:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="60" lane="6" heat="4" heatid="40031" swimtime="00:00:24.31" reactiontime="+63" points="570">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:24.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202730" lastname="BEIQI" firstname="Hana" gender="F" birthdate="2008-09-28">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.83" eventid="13" heat="3" lane="6">
                  <MEETINFO date="2022-07-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.82" eventid="30" heat="3" lane="4">
                  <MEETINFO date="2022-08-15" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="47" lane="6" heat="3" heatid="30013" swimtime="00:00:59.03" reactiontime="+67" points="616">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:28.12" />
                    <SPLIT distance="75" swimtime="00:00:43.70" />
                    <SPLIT distance="100" swimtime="00:00:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="38" lane="4" heat="3" heatid="30030" swimtime="00:00:26.84" reactiontime="+68" points="623">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Saudi Arabia" shortname="KSA" code="KSA" nation="KSA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197181" lastname="ALMAHER" firstname="Mohammed Saeed A" gender="M" birthdate="2007-08-30">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.48" eventid="16" heat="1" lane="3">
                  <MEETINFO date="2021-10-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="29" heat="1" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="58" lane="3" heat="1" heatid="10016" swimtime="00:01:08.84" reactiontime="+65" points="517">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.06" />
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="75" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="-1" lane="3" heat="1" heatid="10029" swimtime="00:02:29.73" status="DSQ" reactiontime="+62" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202026" lastname="ALAYED" firstname="Mashael Meshari A" gender="F" birthdate="2006-12-18">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="13" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="60" lane="4" heat="1" heatid="10013" swimtime="00:01:06.59" reactiontime="+66" points="429">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="75" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:01:06.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="52" lane="6" heat="1" heatid="10030" swimtime="00:00:29.87" reactiontime="+71" points="452">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Kuwait" shortname="KUW" code="KUW" nation="KUW" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="213036" lastname="ZUBAID" firstname="Mohamad" gender="M" birthdate="2008-03-30">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.70" eventid="3" heat="2" lane="1">
                  <MEETINFO date="2022-07-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.30" eventid="14" heat="2" lane="7">
                  <MEETINFO date="2022-07-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="-1" lane="1" heat="2" heatid="20003" swimtime="NT" status="DSQ" />
                <RESULT eventid="14" place="76" lane="7" heat="2" heatid="20014" swimtime="00:00:54.95" reactiontime="+76" points="543">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.69" />
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                    <SPLIT distance="75" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:00:54.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147301" lastname="ALTARMOOM" firstname="Rashed" gender="M" birthdate="1999-04-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.87" eventid="16" heat="2" lane="6">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.35" eventid="41" heat="4" lane="1">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="41" lane="6" heat="2" heatid="20016" swimtime="00:01:00.22" reactiontime="+62" points="773">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="75" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:00.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="37" lane="1" heat="4" heatid="40041" swimtime="00:00:27.66" reactiontime="+62" points="733">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="147305" lastname="DASHTI" firstname="Lara" gender="F" birthdate="2004-01-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.25" eventid="15" heat="2" lane="2">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:35.14" eventid="40" heat="3" lane="7">
                  <MEETINFO date="2021-10-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="47" lane="2" heat="2" heatid="20015" swimtime="00:01:14.61" reactiontime="+68" points="583">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="75" swimtime="00:00:55.07" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="35" lane="7" heat="3" heatid="30040" swimtime="00:00:34.21" reactiontime="+72" points="581">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.00" />
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213037" lastname="SULTAN" firstname="Saba" gender="F" birthdate="2008-05-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.74" eventid="13" heat="2" lane="3">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.20" eventid="30" heat="2" lane="5">
                  <MEETINFO date="2022-07-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="58" lane="3" heat="2" heatid="20013" swimtime="00:01:04.62" reactiontime="+68" points="470">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.58" />
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="75" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="48" lane="5" heat="2" heatid="20030" swimtime="00:00:29.04" reactiontime="+68" points="492">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Latvia" shortname="LAT" code="LAT" nation="LAT" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="130703" lastname="FELDBERGS" firstname="Girts" gender="M" birthdate="1993-02-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.81" eventid="3" heat="3" lane="5">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.62" eventid="19" heat="2" lane="1">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="26" lane="5" heat="3" heatid="30003" swimtime="00:00:52.44" reactiontime="+65" points="782">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:25.12" />
                    <SPLIT distance="75" swimtime="00:00:38.55" />
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="33" lane="1" heat="2" heatid="20019" swimtime="00:00:24.67" reactiontime="+61" points="730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.14" />
                    <SPLIT distance="50" swimtime="00:00:24.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121592" lastname="BOBROVS" firstname="Daniils" gender="M" birthdate="1997-10-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.13" eventid="16" heat="3" lane="4">
                  <MEETINFO date="2021-10-07" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.41" eventid="29" heat="2" lane="5">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="46" lane="4" heat="3" heatid="30016" swimtime="00:01:01.02" reactiontime="+62" points="743">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="75" swimtime="00:00:44.88" />
                    <SPLIT distance="100" swimtime="00:01:01.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="25" lane="5" heat="2" heatid="20029" swimtime="00:02:11.37" reactiontime="+68" points="765">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="75" swimtime="00:00:46.75" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="125" swimtime="00:01:20.66" />
                    <SPLIT distance="150" swimtime="00:01:37.61" />
                    <SPLIT distance="175" swimtime="00:01:54.63" />
                    <SPLIT distance="200" swimtime="00:02:11.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197066" lastname="MIĶELSONS" firstname="Kristaps" gender="M" birthdate="2004-02-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:58.30" eventid="7" heat="2" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:04:15.90" eventid="37" heat="1" lane="3">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="29" lane="5" heat="2" heatid="20007" swimtime="00:01:59.49" reactiontime="+72" points="772">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                    <SPLIT distance="75" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:00:56.27" />
                    <SPLIT distance="125" swimtime="00:01:13.18" />
                    <SPLIT distance="150" swimtime="00:01:30.51" />
                    <SPLIT distance="175" swimtime="00:01:46.15" />
                    <SPLIT distance="200" swimtime="00:01:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="20" lane="3" heat="1" heatid="10037" swimtime="00:04:19.33" reactiontime="+76" points="742">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:27.87" />
                    <SPLIT distance="75" swimtime="00:00:43.93" />
                    <SPLIT distance="100" swimtime="00:01:00.45" />
                    <SPLIT distance="125" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:01:33.66" />
                    <SPLIT distance="175" swimtime="00:01:49.90" />
                    <SPLIT distance="200" swimtime="00:02:05.75" />
                    <SPLIT distance="225" swimtime="00:02:23.83" />
                    <SPLIT distance="250" swimtime="00:02:42.34" />
                    <SPLIT distance="275" swimtime="00:03:00.45" />
                    <SPLIT distance="300" swimtime="00:03:19.01" />
                    <SPLIT distance="325" swimtime="00:03:35.30" />
                    <SPLIT distance="350" swimtime="00:03:50.34" />
                    <SPLIT distance="375" swimtime="00:04:05.21" />
                    <SPLIT distance="400" swimtime="00:04:19.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108263" lastname="BAIKOVA" firstname="Arina" gender="F" birthdate="2000-09-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.44" eventid="13" heat="5" lane="3">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.72" eventid="22" heat="3" lane="8">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="45" lane="3" heat="5" heatid="50013" swimtime="00:00:58.27" reactiontime="+70" points="641">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="75" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:00:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="25" lane="8" heat="3" heatid="30022" swimtime="00:01:05.22" reactiontime="+68" points="650">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:29.08" />
                    <SPLIT distance="75" swimtime="00:00:49.39" />
                    <SPLIT distance="100" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Libya" shortname="LBA" code="LBA" nation="LBA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197567" lastname="ASHOUR" firstname="Abdulhai Abdulmenem Sh" gender="M" birthdate="2006-07-01">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.68" eventid="39" heat="2" lane="6">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="23" heat="2" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="51" lane="6" heat="2" heatid="20039" swimtime="00:01:00.26" reactiontime="+75" points="498">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="75" swimtime="00:00:44.10" />
                    <SPLIT distance="100" swimtime="00:01:00.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="35" lane="8" heat="2" heatid="20023" swimtime="00:01:03.95" reactiontime="+76" points="457">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.79" />
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="75" swimtime="00:00:49.13" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="146394" lastname="QATAT" firstname="Ezuldeen" gender="M" birthdate="1999-05-03">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5" heat="2" lane="3" />
                <ENTRY entrytime="NT" eventid="31" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="65" lane="3" heat="2" heatid="20005" swimtime="00:00:29.48" reactiontime="+76" points="401">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.38" />
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="70" lane="5" heat="1" heatid="10031" swimtime="00:00:26.52" reactiontime="+77" points="439">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Lebanon" shortname="LBN" code="LBN" nation="LBN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="126096" lastname="KHOURY" firstname="Marie" gender="F" birthdate="2001-05-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:28.74" eventid="18" heat="4" lane="7">
                  <MEETINFO date="2021-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.31" eventid="30" heat="4" lane="2">
                  <MEETINFO date="2021-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="37" lane="7" heat="4" heatid="40018" swimtime="00:00:29.35" reactiontime="+54" points="638">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.37" />
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="36" lane="2" heat="4" heatid="40030" swimtime="00:00:26.42" reactiontime="+63" points="653">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:26.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110713" lastname="DOUEIHY" firstname="Gabriella" gender="F" birthdate="1999-04-30">
              <ENTRIES>
                <ENTRY entrytime="00:09:11.65" eventid="12" heat="1" lane="2">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:17:17.12" eventid="33" heat="1" lane="5">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="21" lane="2" heat="1" heatid="10012" swimtime="00:09:11.60" reactiontime="+66" points="656">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="75" swimtime="00:00:47.33" />
                    <SPLIT distance="100" swimtime="00:01:04.19" />
                    <SPLIT distance="125" swimtime="00:01:21.17" />
                    <SPLIT distance="150" swimtime="00:01:38.29" />
                    <SPLIT distance="175" swimtime="00:01:55.56" />
                    <SPLIT distance="200" swimtime="00:02:12.76" />
                    <SPLIT distance="225" swimtime="00:02:30.12" />
                    <SPLIT distance="250" swimtime="00:02:47.50" />
                    <SPLIT distance="275" swimtime="00:03:05.00" />
                    <SPLIT distance="300" swimtime="00:03:22.43" />
                    <SPLIT distance="325" swimtime="00:03:39.94" />
                    <SPLIT distance="350" swimtime="00:03:57.48" />
                    <SPLIT distance="375" swimtime="00:04:15.19" />
                    <SPLIT distance="400" swimtime="00:04:32.74" />
                    <SPLIT distance="425" swimtime="00:04:50.24" />
                    <SPLIT distance="450" swimtime="00:05:07.86" />
                    <SPLIT distance="475" swimtime="00:05:25.42" />
                    <SPLIT distance="500" swimtime="00:05:42.81" />
                    <SPLIT distance="525" swimtime="00:06:00.37" />
                    <SPLIT distance="550" swimtime="00:06:17.98" />
                    <SPLIT distance="575" swimtime="00:06:35.48" />
                    <SPLIT distance="600" swimtime="00:06:53.02" />
                    <SPLIT distance="625" swimtime="00:07:10.63" />
                    <SPLIT distance="650" swimtime="00:07:28.39" />
                    <SPLIT distance="675" swimtime="00:07:45.87" />
                    <SPLIT distance="700" swimtime="00:08:03.48" />
                    <SPLIT distance="725" swimtime="00:08:20.88" />
                    <SPLIT distance="750" swimtime="00:08:38.31" />
                    <SPLIT distance="775" swimtime="00:08:55.26" />
                    <SPLIT distance="800" swimtime="00:09:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="17" lane="5" heat="1" heatid="10033" swimtime="00:17:20.28" reactiontime="+61" points="687">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.42" />
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="75" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:04.04" />
                    <SPLIT distance="125" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:01:38.23" />
                    <SPLIT distance="175" swimtime="00:01:55.57" />
                    <SPLIT distance="200" swimtime="00:02:12.95" />
                    <SPLIT distance="225" swimtime="00:02:30.26" />
                    <SPLIT distance="250" swimtime="00:02:47.34" />
                    <SPLIT distance="275" swimtime="00:03:04.53" />
                    <SPLIT distance="300" swimtime="00:03:21.85" />
                    <SPLIT distance="325" swimtime="00:03:39.07" />
                    <SPLIT distance="350" swimtime="00:03:56.50" />
                    <SPLIT distance="375" swimtime="00:04:13.92" />
                    <SPLIT distance="400" swimtime="00:04:31.12" />
                    <SPLIT distance="425" swimtime="00:04:48.71" />
                    <SPLIT distance="450" swimtime="00:05:05.99" />
                    <SPLIT distance="475" swimtime="00:05:23.55" />
                    <SPLIT distance="500" swimtime="00:05:41.11" />
                    <SPLIT distance="525" swimtime="00:05:58.82" />
                    <SPLIT distance="550" swimtime="00:06:16.23" />
                    <SPLIT distance="575" swimtime="00:06:33.89" />
                    <SPLIT distance="600" swimtime="00:06:51.40" />
                    <SPLIT distance="625" swimtime="00:07:09.00" />
                    <SPLIT distance="650" swimtime="00:07:26.51" />
                    <SPLIT distance="675" swimtime="00:07:44.04" />
                    <SPLIT distance="700" swimtime="00:08:01.43" />
                    <SPLIT distance="725" swimtime="00:08:19.01" />
                    <SPLIT distance="750" swimtime="00:08:36.47" />
                    <SPLIT distance="775" swimtime="00:08:53.91" />
                    <SPLIT distance="800" swimtime="00:09:11.15" />
                    <SPLIT distance="825" swimtime="00:09:28.77" />
                    <SPLIT distance="850" swimtime="00:09:46.46" />
                    <SPLIT distance="875" swimtime="00:10:04.00" />
                    <SPLIT distance="900" swimtime="00:10:21.50" />
                    <SPLIT distance="925" swimtime="00:10:38.96" />
                    <SPLIT distance="950" swimtime="00:10:56.44" />
                    <SPLIT distance="975" swimtime="00:11:14.10" />
                    <SPLIT distance="1000" swimtime="00:11:31.67" />
                    <SPLIT distance="1025" swimtime="00:11:49.26" />
                    <SPLIT distance="1050" swimtime="00:12:06.76" />
                    <SPLIT distance="1075" swimtime="00:12:24.50" />
                    <SPLIT distance="1100" swimtime="00:12:41.87" />
                    <SPLIT distance="1125" swimtime="00:12:59.45" />
                    <SPLIT distance="1150" swimtime="00:13:17.29" />
                    <SPLIT distance="1175" swimtime="00:13:34.74" />
                    <SPLIT distance="1200" swimtime="00:13:52.43" />
                    <SPLIT distance="1225" swimtime="00:14:10.11" />
                    <SPLIT distance="1250" swimtime="00:14:27.67" />
                    <SPLIT distance="1275" swimtime="00:14:45.08" />
                    <SPLIT distance="1300" swimtime="00:15:02.51" />
                    <SPLIT distance="1325" swimtime="00:15:20.06" />
                    <SPLIT distance="1350" swimtime="00:15:37.51" />
                    <SPLIT distance="1375" swimtime="00:15:55.28" />
                    <SPLIT distance="1400" swimtime="00:16:12.60" />
                    <SPLIT distance="1425" swimtime="00:16:29.87" />
                    <SPLIT distance="1450" swimtime="00:16:47.11" />
                    <SPLIT distance="1475" swimtime="00:17:04.25" />
                    <SPLIT distance="1500" swimtime="00:17:20.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Lithuania" shortname="LTU" code="LTU" nation="LTU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="124935" lastname="SIDLAUSKAS" firstname="Andrius" gender="M" birthdate="1997-04-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.52" eventid="16" heat="8" lane="7">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.14" eventid="29" heat="5" lane="2">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.22" eventid="41" heat="9" lane="2">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="30" lane="7" heat="8" heatid="80016" swimtime="00:00:58.60" reactiontime="+65" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="75" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:00:58.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="21" lane="2" heat="5" heatid="50029" swimtime="00:02:08.69" reactiontime="+66" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="75" swimtime="00:00:44.53" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="125" swimtime="00:01:16.81" />
                    <SPLIT distance="150" swimtime="00:01:33.41" />
                    <SPLIT distance="175" swimtime="00:01:50.72" />
                    <SPLIT distance="200" swimtime="00:02:08.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="22" lane="2" heat="9" heatid="90041" swimtime="00:00:26.80" reactiontime="+66" points="806">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101986" lastname="RAPSYS" firstname="Danas" gender="M" birthdate="1995-05-21">
              <ENTRIES>
                <ENTRY entrytime="00:01:41.17" eventid="44" heat="6" lane="5">
                  <MEETINFO date="2021-10-03" />
                </ENTRY>
                <ENTRY entrytime="00:03:36.23" eventid="24" heat="4" lane="4">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="144" place="7" lane="2" heat="1" heatid="10144" swimtime="00:01:41.74" reactiontime="+65" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.21" />
                    <SPLIT distance="50" swimtime="00:00:23.84" />
                    <SPLIT distance="75" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:00:49.66" />
                    <SPLIT distance="125" swimtime="00:01:02.79" />
                    <SPLIT distance="150" swimtime="00:01:15.95" />
                    <SPLIT distance="175" swimtime="00:01:29.00" />
                    <SPLIT distance="200" swimtime="00:01:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="5" lane="5" heat="6" heatid="60044" swimtime="00:01:42.21" reactiontime="+65" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:24.09" />
                    <SPLIT distance="75" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:00:50.49" />
                    <SPLIT distance="125" swimtime="00:01:03.72" />
                    <SPLIT distance="150" swimtime="00:01:16.86" />
                    <SPLIT distance="175" swimtime="00:01:29.71" />
                    <SPLIT distance="200" swimtime="00:01:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="124" place="3" lane="1" heat="1" heatid="10124" swimtime="00:03:36.26" reactiontime="+66" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:25.03" />
                    <SPLIT distance="75" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:00:52.21" />
                    <SPLIT distance="125" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:19.74" />
                    <SPLIT distance="175" swimtime="00:01:33.63" />
                    <SPLIT distance="200" swimtime="00:01:47.44" />
                    <SPLIT distance="225" swimtime="00:02:01.39" />
                    <SPLIT distance="250" swimtime="00:02:15.23" />
                    <SPLIT distance="275" swimtime="00:02:29.09" />
                    <SPLIT distance="300" swimtime="00:02:42.73" />
                    <SPLIT distance="325" swimtime="00:02:56.50" />
                    <SPLIT distance="350" swimtime="00:03:10.10" />
                    <SPLIT distance="375" swimtime="00:03:23.43" />
                    <SPLIT distance="400" swimtime="00:03:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="7" lane="4" heat="4" heatid="40024" swimtime="00:03:38.71" reactiontime="+68" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:25.10" />
                    <SPLIT distance="75" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:00:52.65" />
                    <SPLIT distance="125" swimtime="00:01:06.49" />
                    <SPLIT distance="150" swimtime="00:01:20.45" />
                    <SPLIT distance="175" swimtime="00:01:34.37" />
                    <SPLIT distance="200" swimtime="00:01:48.33" />
                    <SPLIT distance="225" swimtime="00:02:02.31" />
                    <SPLIT distance="250" swimtime="00:02:16.29" />
                    <SPLIT distance="275" swimtime="00:02:30.21" />
                    <SPLIT distance="300" swimtime="00:02:44.21" />
                    <SPLIT distance="325" swimtime="00:02:58.12" />
                    <SPLIT distance="350" swimtime="00:03:12.09" />
                    <SPLIT distance="375" swimtime="00:03:25.59" />
                    <SPLIT distance="400" swimtime="00:03:38.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102069" lastname="MEILUTYTE" firstname="Ruta" gender="F" birthdate="1997-03-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.77" eventid="15" heat="7" lane="4">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.60" eventid="40" heat="7" lane="4">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="-1" lane="5" heat="1" heatid="10115" swimtime="00:01:02.91" status="DSQ" reactiontime="+57" />
                <RESULT eventid="15" place="1" lane="4" heat="7" heatid="70015" swimtime="00:01:03.81" reactiontime="+60" points="933">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.40" />
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="75" swimtime="00:00:46.40" />
                    <SPLIT distance="100" swimtime="00:01:03.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="2" lane="4" heat="2" heatid="20215" swimtime="00:01:03.40" reactiontime="+60" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                    <SPLIT distance="75" swimtime="00:00:46.13" />
                    <SPLIT distance="100" swimtime="00:01:03.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="1" lane="4" heat="1" heatid="10140" swimtime="00:00:28.50" reactiontime="+58" points="1006">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="1" lane="4" heat="7" heatid="70040" swimtime="00:00:29.10" reactiontime="+59" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="1" lane="4" heat="2" heatid="20240" swimtime="00:00:28.37" reactiontime="+58" points="1020">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154270" lastname="TETEREVKOVA" firstname="Kotryna" gender="F" birthdate="2002-01-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.54" eventid="15" heat="7" lane="3">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:20.94" eventid="28" heat="4" lane="6">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.19" eventid="40" heat="7" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="-1" lane="3" heat="7" heatid="70015" swimtime="NT" status="DNS" />
                <RESULT eventid="28" place="-1" lane="6" heat="4" heatid="40028" swimtime="NT" status="DNS" />
                <RESULT eventid="40" place="-1" lane="1" heat="7" heatid="70040" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Luxembourg" shortname="LUX" code="LUX" nation="LUX" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="157504" lastname="MANNES" firstname="Max" gender="M" birthdate="1997-11-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:47.61" eventid="44" heat="2" lane="6">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="24" heat="1" lane="7" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="31" lane="6" heat="2" heatid="20044" swimtime="00:01:47.41" reactiontime="+74" points="791">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:25.14" />
                    <SPLIT distance="75" swimtime="00:00:38.82" />
                    <SPLIT distance="100" swimtime="00:00:52.51" />
                    <SPLIT distance="125" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:19.70" />
                    <SPLIT distance="175" swimtime="00:01:33.77" />
                    <SPLIT distance="200" swimtime="00:01:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="27" lane="7" heat="1" heatid="10024" swimtime="00:03:50.63" reactiontime="+74" points="779">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                    <SPLIT distance="75" swimtime="00:00:40.23" />
                    <SPLIT distance="100" swimtime="00:00:54.40" />
                    <SPLIT distance="125" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:23.21" />
                    <SPLIT distance="175" swimtime="00:01:37.71" />
                    <SPLIT distance="200" swimtime="00:01:52.29" />
                    <SPLIT distance="225" swimtime="00:02:06.71" />
                    <SPLIT distance="250" swimtime="00:02:21.43" />
                    <SPLIT distance="275" swimtime="00:02:36.04" />
                    <SPLIT distance="300" swimtime="00:02:50.84" />
                    <SPLIT distance="325" swimtime="00:03:05.53" />
                    <SPLIT distance="350" swimtime="00:03:20.62" />
                    <SPLIT distance="375" swimtime="00:03:35.82" />
                    <SPLIT distance="400" swimtime="00:03:50.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109083" lastname="HENX" firstname="Julien" gender="M" birthdate="1995-06-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:23.69" eventid="5" heat="5" lane="1">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.08" eventid="31" heat="7" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="38" lane="1" heat="5" heatid="50005" swimtime="00:00:23.30" reactiontime="+63" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.45" />
                    <SPLIT distance="50" swimtime="00:00:23.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="35" lane="1" heat="7" heatid="70031" swimtime="00:00:21.57" reactiontime="+64" points="816">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.29" />
                    <SPLIT distance="50" swimtime="00:00:21.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Sint Maarten" shortname="MAA" code="MAA" nation="MAA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197907" lastname="ILLIS" firstname="Abbi" gender="F" birthdate="2003-12-06">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.97" eventid="13" heat="2" lane="2">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:49.20" eventid="40" heat="2" lane="2">
                  <MEETINFO date="2022-05-15" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="62" lane="2" heat="2" heatid="20013" swimtime="00:01:09.62" reactiontime="+66" points="376">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="75" swimtime="00:00:51.37" />
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="42" lane="2" heat="2" heatid="20040" swimtime="00:00:42.87" reactiontime="+66" points="295">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.18" />
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="167035" lastname="ILLIS" firstname="Taffi" gender="F" birthdate="2001-09-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:31.25" eventid="4" heat="2" lane="6">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.11" eventid="30" heat="3" lane="7">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="36" lane="6" heat="2" heatid="20004" swimtime="00:00:31.16" reactiontime="+61" points="478">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.20" />
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="51" lane="7" heat="3" heatid="30030" swimtime="00:00:29.77" reactiontime="+63" points="456">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Macau, China" shortname="MAC" code="MAC" nation="MAC" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="108152" lastname="CHAO" firstname="Man Hou" gender="M" birthdate="1996-02-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.01" eventid="16" heat="5" lane="4">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.74" eventid="41" heat="8" lane="8">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="18" lane="4" heat="5" heatid="50016" swimtime="00:00:58.01" reactiontime="+69" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                    <SPLIT distance="75" swimtime="00:00:42.42" />
                    <SPLIT distance="100" swimtime="00:00:58.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="14" lane="8" heat="8" heatid="80041" swimtime="00:00:26.46" reactiontime="+68" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="16" lane="1" heat="1" heatid="10241" swimtime="00:00:26.77" reactiontime="+69" points="809">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.27" />
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118815" lastname="LIN" firstname="Sizhuang" gender="M" birthdate="1999-03-29">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="7" heat="1" lane="6" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="42" heat="1" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="34" lane="6" heat="1" heatid="10007" swimtime="00:02:02.41" reactiontime="+70" points="718">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                    <SPLIT distance="75" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:00:57.92" />
                    <SPLIT distance="125" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:01:33.41" />
                    <SPLIT distance="175" swimtime="00:01:48.43" />
                    <SPLIT distance="200" swimtime="00:02:02.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="22" lane="8" heat="1" heatid="10042" swimtime="00:08:21.81" reactiontime="+71" points="689">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.51" />
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="75" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:00:58.63" />
                    <SPLIT distance="125" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:01:29.54" />
                    <SPLIT distance="175" swimtime="00:01:45.16" />
                    <SPLIT distance="200" swimtime="00:02:00.99" />
                    <SPLIT distance="225" swimtime="00:02:16.66" />
                    <SPLIT distance="250" swimtime="00:02:32.58" />
                    <SPLIT distance="275" swimtime="00:02:48.39" />
                    <SPLIT distance="300" swimtime="00:03:04.24" />
                    <SPLIT distance="325" swimtime="00:03:20.06" />
                    <SPLIT distance="350" swimtime="00:03:35.93" />
                    <SPLIT distance="375" swimtime="00:03:51.71" />
                    <SPLIT distance="400" swimtime="00:04:07.54" />
                    <SPLIT distance="425" swimtime="00:04:23.37" />
                    <SPLIT distance="450" swimtime="00:04:39.20" />
                    <SPLIT distance="475" swimtime="00:04:54.87" />
                    <SPLIT distance="500" swimtime="00:05:10.55" />
                    <SPLIT distance="525" swimtime="00:05:26.20" />
                    <SPLIT distance="550" swimtime="00:05:41.87" />
                    <SPLIT distance="575" swimtime="00:05:57.52" />
                    <SPLIT distance="600" swimtime="00:06:13.26" />
                    <SPLIT distance="625" swimtime="00:06:29.06" />
                    <SPLIT distance="650" swimtime="00:06:45.12" />
                    <SPLIT distance="675" swimtime="00:07:01.33" />
                    <SPLIT distance="700" swimtime="00:07:17.70" />
                    <SPLIT distance="725" swimtime="00:07:33.89" />
                    <SPLIT distance="750" swimtime="00:07:50.11" />
                    <SPLIT distance="775" swimtime="00:08:06.18" />
                    <SPLIT distance="800" swimtime="00:08:21.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118818" lastname="CHEANG" firstname="Weng Lam" gender="F" birthdate="2000-11-16">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="2" heat="1" lane="2" />
                <ENTRY entrytime="NT" eventid="18" heat="2" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="40" lane="2" heat="1" heatid="10002" swimtime="00:01:04.74" reactiontime="+64" points="609">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.34" />
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="75" swimtime="00:00:48.30" />
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="41" lane="8" heat="2" heatid="20018" swimtime="00:00:30.24" reactiontime="+61" points="583">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.16" />
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212765" lastname="CHEN" firstname="Pui Lam" gender="F" birthdate="2008-01-08">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="15" heat="1" lane="7" />
                <ENTRY entrytime="NT" eventid="6" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="38" lane="7" heat="1" heatid="10015" swimtime="00:01:09.79" reactiontime="+72" points="713">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="75" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="33" lane="5" heat="1" heatid="10006" swimtime="00:02:23.61" reactiontime="+71" points="610">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="75" swimtime="00:00:49.68" />
                    <SPLIT distance="100" swimtime="00:01:08.69" />
                    <SPLIT distance="125" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:01:48.69" />
                    <SPLIT distance="175" swimtime="00:02:07.25" />
                    <SPLIT distance="200" swimtime="00:02:23.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Macau, China">
              <RESULTS>
                <RESULT eventid="27" place="18" lane="1" heat="3" swimtime="00:01:38.91" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.94" />
                    <SPLIT distance="50" swimtime="00:00:22.60" />
                    <SPLIT distance="75" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:00:45.57" />
                    <SPLIT distance="125" swimtime="00:00:58.46" />
                    <SPLIT distance="150" swimtime="00:01:12.21" />
                    <SPLIT distance="175" swimtime="00:01:25.05" />
                    <SPLIT distance="200" swimtime="00:01:38.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="108152" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="118815" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="118818" reactiontime="+40" />
                    <RELAYPOSITION number="4" athleteid="212765" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Madagascar" shortname="MAD" code="MAD" nation="MAD" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="163157" lastname="RAHARVEL" firstname="Jonathan" gender="M" birthdate="2002-04-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.73" eventid="16" heat="2" lane="5">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.82" eventid="41" heat="3" lane="5">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="50" lane="5" heat="2" heatid="20016" swimtime="00:01:01.84" reactiontime="+63" points="714">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="75" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="47" lane="5" heat="3" heatid="30041" swimtime="00:00:28.55" reactiontime="+63" points="667">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163217" lastname="TENDRINAVALONA" firstname="Idealy" gender="F" birthdate="2004-07-02">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="2" heat="1" lane="1" />
                <ENTRY entrytime="NT" eventid="18" heat="1" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="43" lane="1" heat="1" heatid="10002" swimtime="00:01:08.30" reactiontime="+62" points="519">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.80" />
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="75" swimtime="00:00:50.00" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="42" lane="3" heat="1" heatid="10018" swimtime="00:00:32.19" reactiontime="+58" points="483">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.47" />
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Malawi" shortname="MAW" code="MAW" nation="MAW" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="138512" lastname="GOMES" firstname="Filipe" gender="M" birthdate="1997-04-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.92" eventid="5" heat="3" lane="5">
                  <MEETINFO date="2021-11-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="23" heat="1" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="55" lane="5" heat="3" heatid="30005" swimtime="00:00:25.90" reactiontime="+62" points="592">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="34" lane="6" heat="1" heatid="10023" swimtime="00:00:58.44" reactiontime="+61" points="599">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="75" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:00:58.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="113630" lastname="PINTO" firstname="Ammara" gender="F" birthdate="1997-09-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.60" eventid="13" heat="3" lane="8">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.75" eventid="30" heat="3" lane="1">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="61" lane="8" heat="3" heatid="30013" swimtime="00:01:07.47" reactiontime="+64" points="413">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="75" swimtime="00:00:50.14" />
                    <SPLIT distance="100" swimtime="00:01:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="49" lane="1" heat="3" heatid="30030" swimtime="00:00:29.71" reactiontime="+61" points="459">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.28" />
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161267" lastname="MAKWENDA" firstname="Jessica" gender="F" birthdate="2005-10-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:39.32" eventid="40" heat="2" lane="5">
                  <MEETINFO date="2021-10-13" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.07" eventid="4" heat="2" lane="7">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="39" lane="5" heat="2" heatid="20040" swimtime="00:00:38.99" reactiontime="+72" points="393">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.23" />
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="40" lane="7" heat="2" heatid="20004" swimtime="00:00:35.18" reactiontime="+70" points="332">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Rep. of Moldova" shortname="MDA" code="MDA" nation="MDA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="164543" lastname="MALACHI" firstname="Constantin" gender="M" birthdate="1997-04-11">
              <ENTRIES>
                <ENTRY entrytime="00:02:10.39" eventid="29" heat="2" lane="6">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.52" eventid="41" heat="5" lane="2">
                  <MEETINFO date="2022-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="29" place="-1" lane="6" heat="2" heatid="20029" swimtime="NT" status="DNS" />
                <RESULT eventid="41" place="36" lane="2" heat="5" heatid="50041" swimtime="00:00:27.63" reactiontime="+66" points="736">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196969" lastname="ALOVAȚKI" firstname="Pavel" gender="M" birthdate="2003-10-31">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.26" eventid="44" heat="1" lane="4">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:03:55.64" eventid="24" heat="2" lane="1">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="41" lane="4" heat="1" heatid="10044" swimtime="00:01:51.42" reactiontime="+62" points="709">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                    <SPLIT distance="50" swimtime="00:00:26.61" />
                    <SPLIT distance="75" swimtime="00:00:40.76" />
                    <SPLIT distance="100" swimtime="00:00:55.16" />
                    <SPLIT distance="125" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:23.82" />
                    <SPLIT distance="175" swimtime="00:01:38.07" />
                    <SPLIT distance="200" swimtime="00:01:51.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="30" lane="1" heat="2" heatid="20024" swimtime="00:03:56.60" reactiontime="+63" points="721">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.47" />
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="75" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:00:56.64" />
                    <SPLIT distance="125" swimtime="00:01:11.47" />
                    <SPLIT distance="150" swimtime="00:01:26.45" />
                    <SPLIT distance="175" swimtime="00:01:41.43" />
                    <SPLIT distance="200" swimtime="00:01:56.42" />
                    <SPLIT distance="225" swimtime="00:02:11.28" />
                    <SPLIT distance="250" swimtime="00:02:26.37" />
                    <SPLIT distance="275" swimtime="00:02:41.57" />
                    <SPLIT distance="300" swimtime="00:02:56.75" />
                    <SPLIT distance="325" swimtime="00:03:11.88" />
                    <SPLIT distance="350" swimtime="00:03:27.00" />
                    <SPLIT distance="375" swimtime="00:03:42.25" />
                    <SPLIT distance="400" swimtime="00:03:56.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="128891" lastname="SALCUTAN" firstname="Tatiana" gender="F" birthdate="2001-04-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.73" eventid="2" heat="2" lane="5">
                  <MEETINFO date="2022-05-15" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.45" eventid="45" heat="2" lane="2">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="34" lane="5" heat="2" heatid="20002" swimtime="00:01:01.16" reactiontime="+68" points="722">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="75" swimtime="00:00:45.17" />
                    <SPLIT distance="100" swimtime="00:01:01.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="-1" lane="2" heat="2" heatid="20045" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Maldives" shortname="MDV" code="MDV" nation="MDV" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="211066" lastname="SHIHAM" firstname="Mohamed Rihan" gender="M" birthdate="2006-12-31">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.87" eventid="3" heat="1" lane="5">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:34.77" eventid="21" heat="1" lane="5">
                  <MEETINFO date="2022-09-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="40" lane="5" heat="1" heatid="10003" swimtime="00:01:07.35" reactiontime="+76" points="369">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="75" swimtime="00:00:50.35" />
                    <SPLIT distance="100" swimtime="00:01:07.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="27" lane="5" heat="1" heatid="10021" swimtime="00:02:27.12" reactiontime="+79" points="398">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="75" swimtime="00:00:50.59" />
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                    <SPLIT distance="125" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                    <SPLIT distance="175" swimtime="00:02:08.80" />
                    <SPLIT distance="200" swimtime="00:02:27.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109057" lastname="IBRAHIM" firstname="Mubal Azzam" gender="M" birthdate="2000-11-03">
              <ENTRIES>
                <ENTRY entrytime="00:02:23.69" eventid="7" heat="1" lane="3">
                  <MEETINFO date="2022-08-03" />
                </ENTRY>
                <ENTRY entrytime="00:05:14.91" eventid="37" heat="1" lane="1">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="36" lane="3" heat="1" heatid="10007" swimtime="00:02:19.77" reactiontime="+65" points="482">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:48.80" />
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                    <SPLIT distance="125" swimtime="00:01:27.15" />
                    <SPLIT distance="150" swimtime="00:01:48.06" />
                    <SPLIT distance="175" swimtime="00:02:04.60" />
                    <SPLIT distance="200" swimtime="00:02:19.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="21" lane="1" heat="1" heatid="10037" swimtime="00:05:00.64" reactiontime="+63" points="476">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="75" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:06.97" />
                    <SPLIT distance="125" swimtime="00:01:27.04" />
                    <SPLIT distance="150" swimtime="00:01:46.65" />
                    <SPLIT distance="175" swimtime="00:02:06.01" />
                    <SPLIT distance="200" swimtime="00:02:25.18" />
                    <SPLIT distance="225" swimtime="00:02:46.83" />
                    <SPLIT distance="250" swimtime="00:03:08.46" />
                    <SPLIT distance="275" swimtime="00:03:30.32" />
                    <SPLIT distance="300" swimtime="00:03:52.40" />
                    <SPLIT distance="325" swimtime="00:04:09.77" />
                    <SPLIT distance="350" swimtime="00:04:26.64" />
                    <SPLIT distance="375" swimtime="00:04:43.83" />
                    <SPLIT distance="400" swimtime="00:05:00.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130525" lastname="SAUSAN" firstname="Aishath" gender="F" birthdate="1988-06-20">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:14.03" eventid="2" heat="1" lane="3" />
                <ENTRY entrytime="00:00:34.76" eventid="18" heat="2" lane="2">
                  <MEETINFO date="2022-08-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="45" lane="3" heat="1" heatid="10002" swimtime="00:01:14.05" reactiontime="+68" points="407">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.80" />
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="75" swimtime="00:00:54.19" />
                    <SPLIT distance="100" swimtime="00:01:14.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="45" lane="2" heat="2" heatid="20018" swimtime="00:00:33.10" reactiontime="+65" points="444">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.34" />
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156129" lastname="AHMED" firstname="Hamna" gender="F" birthdate="2003-04-18">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="45" heat="1" lane="6" />
                <ENTRY entrytime="00:00:30.61" eventid="30" heat="2" lane="3">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="35" lane="6" heat="1" heatid="10045" swimtime="00:02:59.77" reactiontime="+62" points="289">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.67" />
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="75" swimtime="00:01:01.45" />
                    <SPLIT distance="100" swimtime="00:01:24.62" />
                    <SPLIT distance="125" swimtime="00:01:48.51" />
                    <SPLIT distance="150" swimtime="00:02:12.72" />
                    <SPLIT distance="175" swimtime="00:02:36.71" />
                    <SPLIT distance="200" swimtime="00:02:59.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="54" lane="3" heat="2" heatid="20030" swimtime="00:00:30.35" reactiontime="+66" points="431">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.53" />
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Maldives">
              <RESULTS>
                <RESULT eventid="27" place="26" lane="2" heat="2" swimtime="00:01:52.92" reactiontime="+73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:26.14" />
                    <SPLIT distance="75" swimtime="00:00:40.60" />
                    <SPLIT distance="100" swimtime="00:00:56.06" />
                    <SPLIT distance="125" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:26.94" />
                    <SPLIT distance="175" swimtime="00:01:39.34" />
                    <SPLIT distance="200" swimtime="00:01:52.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109057" reactiontime="+73" />
                    <RELAYPOSITION number="2" athleteid="130525" reactiontime="+46" />
                    <RELAYPOSITION number="3" athleteid="156129" reactiontime="+62" />
                    <RELAYPOSITION number="4" athleteid="211066" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Maldives">
              <RESULTS>
                <RESULT eventid="11" place="31" lane="2" heat="4" swimtime="00:02:05.53" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="75" swimtime="00:00:51.23" />
                    <SPLIT distance="100" swimtime="00:01:11.86" />
                    <SPLIT distance="125" swimtime="00:01:24.78" />
                    <SPLIT distance="150" swimtime="00:01:39.81" />
                    <SPLIT distance="175" swimtime="00:01:52.16" />
                    <SPLIT distance="200" swimtime="00:02:05.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130525" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="156129" reactiontime="+64" />
                    <RELAYPOSITION number="3" athleteid="211066" reactiontime="+60" />
                    <RELAYPOSITION number="4" athleteid="109057" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Mexico" shortname="MEX" code="MEX" nation="MEX" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="124974" lastname="MARTINEZ" firstname="Jose" gender="M" birthdate="1997-06-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.46" eventid="39" heat="6" lane="1">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.58" eventid="21" heat="2" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.72" eventid="5" heat="10" lane="8">
                  <MEETINFO date="2021-11-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="19" lane="1" heat="6" heatid="60039" swimtime="00:00:51.06" reactiontime="+63" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.94" />
                    <SPLIT distance="50" swimtime="00:00:23.68" />
                    <SPLIT distance="75" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:00:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="16" lane="6" heat="2" heatid="20021" swimtime="00:01:53.16" reactiontime="+64" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:25.30" />
                    <SPLIT distance="75" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:00:54.33" />
                    <SPLIT distance="125" swimtime="00:01:08.90" />
                    <SPLIT distance="150" swimtime="00:01:23.71" />
                    <SPLIT distance="175" swimtime="00:01:38.24" />
                    <SPLIT distance="200" swimtime="00:01:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="40" lane="8" heat="10" heatid="100005" swimtime="00:00:23.32" reactiontime="+64" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.71" />
                    <SPLIT distance="50" swimtime="00:00:23.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213739" lastname="GRANA PEREZ" firstname="Miranda" gender="F" birthdate="2004-11-05">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.35" eventid="2" heat="2" lane="6">
                  <MEETINFO date="2022-04-08" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.96" eventid="18" heat="3" lane="6">
                  <MEETINFO date="2022-04-09" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="26" lane="6" heat="2" heatid="20002" swimtime="00:00:58.80" reactiontime="+55" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                    <SPLIT distance="50" swimtime="00:00:28.01" />
                    <SPLIT distance="75" swimtime="00:00:43.26" />
                    <SPLIT distance="100" swimtime="00:00:58.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="24" lane="6" heat="3" heatid="30018" swimtime="00:00:27.17" reactiontime="+51" points="804">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Mongolia" shortname="MGL" code="MGL" nation="MGL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="156544" lastname="BATBAYAR" firstname="Enkhtamir" gender="M" birthdate="2004-09-27">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="39" heat="1" lane="5" />
                <ENTRY entrytime="00:00:52.09" eventid="14" heat="4" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="48" lane="5" heat="1" heatid="10039" swimtime="00:00:57.02" reactiontime="+69" points="588">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:26.27" />
                    <SPLIT distance="75" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:00:57.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="58" lane="2" heat="4" heatid="40014" swimtime="00:00:50.87" reactiontime="+75" points="684">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:24.50" />
                    <SPLIT distance="75" swimtime="00:00:37.82" />
                    <SPLIT distance="100" swimtime="00:00:50.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119363" lastname="MYAGMAR" firstname="Delgerkhuu" gender="M" birthdate="1996-09-21">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="41" heat="1" lane="4" />
                <ENTRY entrytime="00:00:24.63" eventid="31" heat="4" lane="2">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="51" lane="4" heat="1" heatid="10041" swimtime="00:00:29.85" reactiontime="+65" points="583">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="58" lane="2" heat="4" heatid="40031" swimtime="00:00:24.21" reactiontime="+67" points="577">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162409" lastname="ENKH-AMGALAN" firstname="Ariuntamir" gender="F" birthdate="2004-04-08">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:10.31" eventid="2" heat="1" lane="5" />
                <ENTRY entrytime="00:00:31.95" eventid="18" heat="2" lane="4" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="41" lane="5" heat="1" heatid="10002" swimtime="00:01:04.98" reactiontime="+65" points="602">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                    <SPLIT distance="75" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="38" lane="4" heat="2" heatid="20018" swimtime="00:00:29.68" reactiontime="+65" points="617">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.44" />
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119676" lastname="BATBAYAR" firstname="Enkhkhuslen" gender="F" birthdate="2001-12-14">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:56.08" eventid="13" heat="5" lane="1">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:01:58.23" eventid="43" heat="5" lane="8">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="38" lane="1" heat="5" heatid="50013" swimtime="00:00:55.76" reactiontime="+71" points="731">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="75" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:00:55.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="15" lane="8" heat="5" heatid="50043" swimtime="00:01:56.46" reactiontime="+71" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:27.28" />
                    <SPLIT distance="75" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:00:56.17" />
                    <SPLIT distance="125" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:25.86" />
                    <SPLIT distance="175" swimtime="00:01:41.13" />
                    <SPLIT distance="200" swimtime="00:01:56.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Mongolia">
              <RESULTS>
                <RESULT eventid="27" place="20" lane="6" heat="2" swimtime="00:01:40.46" reactiontime="+74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:23.54" />
                    <SPLIT distance="75" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:00:47.35" />
                    <SPLIT distance="125" swimtime="00:00:59.60" />
                    <SPLIT distance="150" swimtime="00:01:13.18" />
                    <SPLIT distance="175" swimtime="00:01:26.08" />
                    <SPLIT distance="200" swimtime="00:01:40.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156544" reactiontime="+74" />
                    <RELAYPOSITION number="2" athleteid="119363" reactiontime="+36" />
                    <RELAYPOSITION number="3" athleteid="119676" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="162409" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Mongolia">
              <RESULTS>
                <RESULT eventid="11" place="24" lane="6" heat="2" swimtime="00:01:49.97" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="75" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:00:58.91" />
                    <SPLIT distance="125" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:24.33" />
                    <SPLIT distance="175" swimtime="00:01:36.51" />
                    <SPLIT distance="200" swimtime="00:01:49.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="162409" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="119363" reactiontime="+5" />
                    <RELAYPOSITION number="3" athleteid="156544" reactiontime="+46" />
                    <RELAYPOSITION number="4" athleteid="119676" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Marshall Islands" shortname="MHL" code="MHL" nation="MHL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="145216" lastname="KINONO" firstname="Phillip" gender="M" birthdate="1997-12-10">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.19" eventid="14" heat="1" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.54" eventid="31" heat="3" lane="1">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="83" lane="5" heat="1" heatid="10014" swimtime="00:01:01.29" reactiontime="+66" points="391">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                    <SPLIT distance="75" swimtime="00:00:44.67" />
                    <SPLIT distance="100" swimtime="00:01:01.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="73" lane="1" heat="3" heatid="30031" swimtime="00:00:26.86" reactiontime="+65" points="422">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="141672" lastname="HEPLER" firstname="Kayla" gender="F" birthdate="2002-03-22">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="18" heat="2" lane="7" />
                <ENTRY entrytime="00:00:30.03" eventid="30" heat="3" lane="8">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="48" lane="7" heat="2" heatid="20018" swimtime="00:00:33.99" reactiontime="+72" points="410">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.68" />
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="53" lane="8" heat="3" heatid="30030" swimtime="00:00:30.31" reactiontime="+62" points="432">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Mali" shortname="MLI" code="MLI" nation="MLI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="128725" lastname="KOUMA" firstname="Sebastien" gender="M" birthdate="1997-04-27">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="16" heat="1" lane="2" />
                <ENTRY entrytime="NT" eventid="41" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="53" lane="2" heat="1" heatid="10016" swimtime="00:01:04.39" reactiontime="+70" points="632">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="75" swimtime="00:00:46.73" />
                    <SPLIT distance="100" swimtime="00:01:04.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="48" lane="5" heat="1" heatid="10041" swimtime="00:00:28.73" reactiontime="+67" points="654">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212965" lastname="TOURE" firstname="Batourou" gender="F" birthdate="1994-06-06">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="15" heat="1" lane="2" />
                <ENTRY entrytime="NT" eventid="40" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="51" lane="2" heat="1" heatid="10015" swimtime="00:01:49.99" reactiontime="+77" points="182">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.29" />
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                    <SPLIT distance="75" swimtime="00:01:19.95" />
                    <SPLIT distance="100" swimtime="00:01:49.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="45" lane="5" heat="1" heatid="10040" swimtime="00:00:48.96" reactiontime="+85" points="198">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.29" />
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Malta" shortname="MLT" code="MLT" nation="MLT" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="182748" lastname="CACHIA" firstname="Dylan" gender="M" birthdate="2001-09-15">
              <ENTRIES>
                <ENTRY entrytime="00:03:57.26" eventid="24" heat="1" lane="5">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:08:11.85" eventid="42" heat="1" lane="2">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="24" place="32" lane="5" heat="1" heatid="10024" swimtime="00:04:05.61" reactiontime="+69" points="645">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:26.72" />
                    <SPLIT distance="75" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:00:55.86" />
                    <SPLIT distance="125" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:26.60" />
                    <SPLIT distance="175" swimtime="00:01:42.18" />
                    <SPLIT distance="200" swimtime="00:01:57.84" />
                    <SPLIT distance="225" swimtime="00:02:13.74" />
                    <SPLIT distance="250" swimtime="00:02:29.80" />
                    <SPLIT distance="275" swimtime="00:02:45.93" />
                    <SPLIT distance="300" swimtime="00:03:02.22" />
                    <SPLIT distance="325" swimtime="00:03:18.38" />
                    <SPLIT distance="350" swimtime="00:03:34.66" />
                    <SPLIT distance="375" swimtime="00:03:50.75" />
                    <SPLIT distance="400" swimtime="00:04:05.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="23" lane="2" heat="1" heatid="10042" swimtime="00:08:22.71" reactiontime="+72" points="686">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:43.03" />
                    <SPLIT distance="100" swimtime="00:00:58.45" />
                    <SPLIT distance="125" swimtime="00:01:14.17" />
                    <SPLIT distance="150" swimtime="00:01:29.80" />
                    <SPLIT distance="175" swimtime="00:01:45.47" />
                    <SPLIT distance="200" swimtime="00:02:01.22" />
                    <SPLIT distance="225" swimtime="00:02:17.11" />
                    <SPLIT distance="250" swimtime="00:02:32.80" />
                    <SPLIT distance="275" swimtime="00:02:48.62" />
                    <SPLIT distance="300" swimtime="00:03:04.42" />
                    <SPLIT distance="325" swimtime="00:03:20.51" />
                    <SPLIT distance="350" swimtime="00:03:36.50" />
                    <SPLIT distance="375" swimtime="00:03:52.58" />
                    <SPLIT distance="400" swimtime="00:04:08.69" />
                    <SPLIT distance="425" swimtime="00:04:24.77" />
                    <SPLIT distance="450" swimtime="00:04:40.71" />
                    <SPLIT distance="475" swimtime="00:04:56.69" />
                    <SPLIT distance="500" swimtime="00:05:12.58" />
                    <SPLIT distance="525" swimtime="00:05:28.36" />
                    <SPLIT distance="550" swimtime="00:05:44.39" />
                    <SPLIT distance="575" swimtime="00:06:00.54" />
                    <SPLIT distance="600" swimtime="00:06:16.52" />
                    <SPLIT distance="625" swimtime="00:06:32.45" />
                    <SPLIT distance="650" swimtime="00:06:48.67" />
                    <SPLIT distance="675" swimtime="00:07:04.69" />
                    <SPLIT distance="700" swimtime="00:07:20.92" />
                    <SPLIT distance="725" swimtime="00:07:36.80" />
                    <SPLIT distance="750" swimtime="00:07:52.80" />
                    <SPLIT distance="775" swimtime="00:08:08.43" />
                    <SPLIT distance="800" swimtime="00:08:22.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182752" lastname="GATT" firstname="Sasha" gender="F" birthdate="2005-06-22">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.69" eventid="43" heat="2" lane="1">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:08:38.74" eventid="12" heat="1" lane="4">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="27" lane="1" heat="2" heatid="20043" swimtime="00:02:03.72" reactiontime="+70" points="708">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="75" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="125" swimtime="00:01:15.69" />
                    <SPLIT distance="150" swimtime="00:01:31.81" />
                    <SPLIT distance="175" swimtime="00:01:48.09" />
                    <SPLIT distance="200" swimtime="00:02:03.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="16" lane="4" heat="1" heatid="10012" swimtime="00:08:40.76" reactiontime="+69" points="779">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="75" swimtime="00:00:46.17" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="125" swimtime="00:01:18.69" />
                    <SPLIT distance="150" swimtime="00:01:35.07" />
                    <SPLIT distance="175" swimtime="00:01:51.51" />
                    <SPLIT distance="200" swimtime="00:02:07.82" />
                    <SPLIT distance="225" swimtime="00:02:24.11" />
                    <SPLIT distance="250" swimtime="00:02:40.55" />
                    <SPLIT distance="275" swimtime="00:02:56.94" />
                    <SPLIT distance="300" swimtime="00:03:13.42" />
                    <SPLIT distance="325" swimtime="00:03:29.79" />
                    <SPLIT distance="350" swimtime="00:03:46.30" />
                    <SPLIT distance="375" swimtime="00:04:02.61" />
                    <SPLIT distance="400" swimtime="00:04:19.07" />
                    <SPLIT distance="425" swimtime="00:04:35.44" />
                    <SPLIT distance="450" swimtime="00:04:51.83" />
                    <SPLIT distance="475" swimtime="00:05:08.19" />
                    <SPLIT distance="500" swimtime="00:05:24.64" />
                    <SPLIT distance="525" swimtime="00:05:41.02" />
                    <SPLIT distance="550" swimtime="00:05:57.24" />
                    <SPLIT distance="575" swimtime="00:06:13.84" />
                    <SPLIT distance="600" swimtime="00:06:30.34" />
                    <SPLIT distance="625" swimtime="00:06:46.97" />
                    <SPLIT distance="650" swimtime="00:07:03.49" />
                    <SPLIT distance="675" swimtime="00:07:20.22" />
                    <SPLIT distance="700" swimtime="00:07:36.73" />
                    <SPLIT distance="725" swimtime="00:07:53.04" />
                    <SPLIT distance="750" swimtime="00:08:09.72" />
                    <SPLIT distance="775" swimtime="00:08:25.54" />
                    <SPLIT distance="800" swimtime="00:08:40.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Mozambique" shortname="MOZ" code="MOZ" nation="MOZ" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197954" lastname="LAWRENCE" firstname="Matthew" gender="M" birthdate="2003-12-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.10" eventid="41" heat="3" lane="3">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.93" eventid="5" heat="4" lane="1">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="-1" lane="3" heat="3" heatid="30041" swimtime="NT" status="DNS" />
                <RESULT eventid="5" place="-1" lane="1" heat="4" heatid="40005" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Mauritius" shortname="MRI" code="MRI" nation="MRI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="102145" lastname="VINCENT" firstname="Bradley" gender="M" birthdate="1991-11-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.29" eventid="14" heat="5" lane="7">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.34" eventid="31" heat="5" lane="7">
                  <MEETINFO date="2022-08-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="-1" lane="7" heat="5" heatid="50014" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="50" lane="7" heat="5" heatid="50031" swimtime="00:00:22.76" reactiontime="+69" points="694">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.87" />
                    <SPLIT distance="50" swimtime="00:00:22.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210414" lastname="TEELUCK" firstname="Anishta" gender="F" birthdate="2001-05-07">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.59" eventid="2" heat="2" lane="7">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.01" eventid="45" heat="1" lane="5">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="39" lane="7" heat="2" heatid="20002" swimtime="00:01:03.44" reactiontime="+57" points="647">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.72" />
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                    <SPLIT distance="75" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:03.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="33" lane="5" heat="1" heatid="10045" swimtime="00:02:13.71" reactiontime="+55" points="703">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.48" />
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="75" swimtime="00:00:48.30" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="125" swimtime="00:01:21.64" />
                    <SPLIT distance="150" swimtime="00:01:38.61" />
                    <SPLIT distance="175" swimtime="00:01:56.02" />
                    <SPLIT distance="200" swimtime="00:02:13.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Namibia" shortname="NAM" code="NAM" nation="NAM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="145974" lastname="WANTENAAR" firstname="Ronan" gender="M" birthdate="2001-02-10">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.35" eventid="16" heat="3" lane="7">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.89" eventid="41" heat="4" lane="4">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="42" lane="7" heat="3" heatid="30016" swimtime="00:01:00.35" reactiontime="+64" points="768">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                    <SPLIT distance="75" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:01:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="35" lane="4" heat="4" heatid="40041" swimtime="00:00:27.45" reactiontime="+58" points="750">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="119425" lastname="SKINNER" firstname="Xander" gender="M" birthdate="1998-03-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.40" eventid="14" heat="7" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.19" eventid="31" heat="6" lane="5">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="44" lane="2" heat="7" heatid="70014" swimtime="00:00:48.45" reactiontime="+66" points="792">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.97" />
                    <SPLIT distance="50" swimtime="00:00:23.09" />
                    <SPLIT distance="75" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:00:48.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="43" lane="5" heat="6" heatid="60031" swimtime="00:00:21.85" reactiontime="+64" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.55" />
                    <SPLIT distance="50" swimtime="00:00:21.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Netherlands" shortname="NED" code="NED" nation="NED" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154353" lastname="CORBEAU" firstname="Caspar" gender="M" birthdate="2001-04-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.33" eventid="16" heat="8" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.17" eventid="29" heat="4" lane="3">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:26.15" eventid="41" heat="9" lane="6">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="10" lane="2" heat="8" heatid="80016" swimtime="00:00:57.53" reactiontime="+68" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.16" />
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                    <SPLIT distance="75" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:00:57.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="13" lane="2" heat="1" heatid="10216" swimtime="00:00:57.73" reactiontime="+68" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.17" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:00:57.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="11" lane="3" heat="4" heatid="40029" swimtime="00:02:05.14" reactiontime="+66" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="75" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:00:59.81" />
                    <SPLIT distance="125" swimtime="00:01:16.08" />
                    <SPLIT distance="150" swimtime="00:01:32.17" />
                    <SPLIT distance="175" swimtime="00:01:48.50" />
                    <SPLIT distance="200" swimtime="00:02:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="23" lane="6" heat="9" heatid="90041" swimtime="00:00:26.83" reactiontime="+65" points="804">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.03" />
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106982" lastname="KORSTANJE" firstname="Nyls" gender="M" birthdate="1999-02-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.49" eventid="39" heat="7" lane="5">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.25" eventid="5" heat="9" lane="3">
                  <MEETINFO date="2022-07-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="15" lane="5" heat="7" heatid="70039" swimtime="00:00:50.59" reactiontime="+63" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.48" />
                    <SPLIT distance="50" swimtime="00:00:23.28" />
                    <SPLIT distance="75" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:00:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="14" lane="8" heat="2" heatid="20239" swimtime="00:00:50.59" reactiontime="+65" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.54" />
                    <SPLIT distance="50" swimtime="00:00:23.37" />
                    <SPLIT distance="75" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:00:50.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="16" lane="3" heat="9" heatid="90005" swimtime="00:00:22.53" reactiontime="+61" points="899">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:22.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="305" place="17" lane="5" heat="1" heatid="10305" swimtime="00:00:22.35" reactiontime="+63" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.06" />
                    <SPLIT distance="50" swimtime="00:00:22.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109044" lastname="PIJNENBURG" firstname="Stan" gender="M" birthdate="1996-11-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.38" eventid="14" heat="11" lane="3">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="32" lane="3" heat="11" heatid="110014" swimtime="00:00:47.56" reactiontime="+65" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.62" />
                    <SPLIT distance="50" swimtime="00:00:22.59" />
                    <SPLIT distance="75" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:00:47.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154356" lastname="KROON" firstname="Luc" gender="M" birthdate="2001-08-30">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.20" eventid="44" heat="6" lane="6">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:03:38.33" eventid="24" heat="5" lane="2">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="00:07:44.35" eventid="42">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="18" lane="6" heat="6" heatid="60044" swimtime="00:01:43.86" reactiontime="+71" points="875">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:24.60" />
                    <SPLIT distance="75" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:00:50.86" />
                    <SPLIT distance="125" swimtime="00:01:03.99" />
                    <SPLIT distance="150" swimtime="00:01:17.30" />
                    <SPLIT distance="175" swimtime="00:01:30.57" />
                    <SPLIT distance="200" swimtime="00:01:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="17" lane="2" heat="5" heatid="50024" swimtime="00:03:44.76" reactiontime="+70" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:25.88" />
                    <SPLIT distance="75" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:00:53.99" />
                    <SPLIT distance="125" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:21.98" />
                    <SPLIT distance="175" swimtime="00:01:36.07" />
                    <SPLIT distance="200" swimtime="00:01:50.05" />
                    <SPLIT distance="225" swimtime="00:02:03.70" />
                    <SPLIT distance="250" swimtime="00:02:17.72" />
                    <SPLIT distance="275" swimtime="00:02:31.88" />
                    <SPLIT distance="300" swimtime="00:02:46.32" />
                    <SPLIT distance="325" swimtime="00:03:00.91" />
                    <SPLIT distance="350" swimtime="00:03:15.63" />
                    <SPLIT distance="375" swimtime="00:03:30.42" />
                    <SPLIT distance="400" swimtime="00:03:44.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154915" lastname="JANSEN" firstname="Thomas" gender="M" birthdate="2001-06-06">
              <ENTRIES>
                <ENTRY entrytime="00:04:07.88" eventid="37" heat="2" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="37" place="11" lane="7" heat="2" heatid="20037" swimtime="00:04:08.29" reactiontime="+71" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="75" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:00:56.76" />
                    <SPLIT distance="125" swimtime="00:01:12.27" />
                    <SPLIT distance="150" swimtime="00:01:27.41" />
                    <SPLIT distance="175" swimtime="00:01:42.67" />
                    <SPLIT distance="200" swimtime="00:01:57.79" />
                    <SPLIT distance="225" swimtime="00:02:15.51" />
                    <SPLIT distance="250" swimtime="00:02:33.20" />
                    <SPLIT distance="275" swimtime="00:02:51.23" />
                    <SPLIT distance="300" swimtime="00:03:09.58" />
                    <SPLIT distance="325" swimtime="00:03:24.77" />
                    <SPLIT distance="350" swimtime="00:03:39.36" />
                    <SPLIT distance="375" swimtime="00:03:53.91" />
                    <SPLIT distance="400" swimtime="00:04:08.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129673" lastname="DE BOER" firstname="Thom" gender="M" birthdate="1991-12-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:20.78" eventid="31" heat="10" lane="5">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="21" lane="5" heat="10" heatid="100031" swimtime="00:00:21.35" reactiontime="+64" points="841">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.16" />
                    <SPLIT distance="50" swimtime="00:00:21.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154357" lastname="SIMONS" firstname="Kenzo" gender="M" birthdate="2001-04-13">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.10" eventid="31" heat="9" lane="3">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="18" lane="3" heat="9" heatid="90031" swimtime="00:00:21.33" reactiontime="+59" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="331" place="18" lane="5" heat="1" heatid="10331" swimtime="00:00:21.28" reactiontime="+60" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:21.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109025" lastname="TOUSSAINT" firstname="Kira" gender="F" birthdate="1994-05-22">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.42" eventid="2" heat="4" lane="4">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.26" eventid="45" heat="4" lane="4">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.73" eventid="18" heat="5" lane="4">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="7" lane="8" heat="1" heatid="10102" swimtime="00:00:56.41" reactiontime="+54" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.22" />
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                    <SPLIT distance="75" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:00:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="5" lane="4" heat="4" heatid="40002" swimtime="00:00:56.62" reactiontime="+54" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                    <SPLIT distance="75" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="8" lane="3" heat="2" heatid="20202" swimtime="00:00:56.54" reactiontime="+54" points="914">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:26.99" />
                    <SPLIT distance="75" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:00:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="8" lane="1" heat="1" heatid="10145" swimtime="00:02:05.20" reactiontime="+59" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.00" />
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="75" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="125" swimtime="00:01:17.05" />
                    <SPLIT distance="150" swimtime="00:01:33.01" />
                    <SPLIT distance="175" swimtime="00:01:49.10" />
                    <SPLIT distance="200" swimtime="00:02:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="7" lane="4" heat="4" heatid="40045" swimtime="00:02:03.40" reactiontime="+59" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.92" />
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                    <SPLIT distance="75" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:00.12" />
                    <SPLIT distance="125" swimtime="00:01:15.76" />
                    <SPLIT distance="150" swimtime="00:01:31.40" />
                    <SPLIT distance="175" swimtime="00:01:47.41" />
                    <SPLIT distance="200" swimtime="00:02:03.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="7" lane="4" heat="5" heatid="50018" swimtime="00:00:26.09" reactiontime="+54" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.97" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="10" lane="6" heat="2" heatid="20218" swimtime="00:00:26.17" reactiontime="+55" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:26.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109026" lastname="DE WAARD" firstname="Maaike" gender="F" birthdate="1996-10-11">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:55.86" eventid="2" heat="4" lane="5">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.95" eventid="38" heat="2" lane="6">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.97" eventid="18" heat="5" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.97" eventid="4" heat="4" lane="5">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="10" lane="5" heat="4" heatid="40002" swimtime="00:00:57.01" reactiontime="+62" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                    <SPLIT distance="75" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:00:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="10" lane="2" heat="1" heatid="10202" swimtime="00:00:56.78" reactiontime="+66" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                    <SPLIT distance="75" swimtime="00:00:41.75" />
                    <SPLIT distance="100" swimtime="00:00:56.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="138" place="7" lane="7" heat="1" heatid="10138" swimtime="00:00:56.52" reactiontime="+72" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.67" />
                    <SPLIT distance="50" swimtime="00:00:25.94" />
                    <SPLIT distance="75" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:00:56.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="6" lane="6" heat="2" heatid="20038" swimtime="00:00:56.67" reactiontime="+75" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                    <SPLIT distance="75" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:00:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="7" lane="3" heat="1" heatid="10238" swimtime="00:00:56.40" reactiontime="+74" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                    <SPLIT distance="75" swimtime="00:00:41.02" />
                    <SPLIT distance="100" swimtime="00:00:56.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="8" lane="8" heat="1" heatid="10118" swimtime="00:00:26.16" reactiontime="+63" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.76" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="11" lane="5" heat="5" heatid="50018" swimtime="00:00:26.32" reactiontime="+62" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:26.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="7" lane="7" heat="2" heatid="20218" swimtime="00:00:26.02" reactiontime="+63" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="104" place="7" lane="6" heat="1" heatid="10104" swimtime="00:00:24.98" reactiontime="+70" points="929">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:24.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="10" lane="5" heat="4" heatid="40004" swimtime="00:00:25.40" reactiontime="+74" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:25.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="4" lane="2" heat="1" heatid="10204" swimtime="00:00:24.92" reactiontime="+70" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.46" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129677" lastname="SCHOUTEN" firstname="Tes" gender="F" birthdate="2000-12-31">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.71" eventid="15" heat="5" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.55" eventid="28" heat="5" lane="5">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="2" lane="6" heat="1" heatid="10115" swimtime="00:01:03.90" reactiontime="+64" points="929">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.80" />
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="75" swimtime="00:00:46.72" />
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="5" lane="3" heat="5" heatid="50015" swimtime="00:01:04.22" reactiontime="+65" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="75" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:04.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="4" lane="3" heat="2" heatid="20215" swimtime="00:01:04.31" reactiontime="+66" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:30.27" />
                    <SPLIT distance="75" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="128" place="3" lane="3" heat="1" heatid="10128" swimtime="00:02:18.19" reactiontime="+67" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="75" swimtime="00:00:48.01" />
                    <SPLIT distance="100" swimtime="00:01:05.70" />
                    <SPLIT distance="125" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:01:41.56" />
                    <SPLIT distance="175" swimtime="00:01:59.47" />
                    <SPLIT distance="200" swimtime="00:02:18.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="3" lane="5" heat="5" heatid="50028" swimtime="00:02:18.70" reactiontime="+65" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.26" />
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="75" swimtime="00:00:48.43" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="125" swimtime="00:01:24.33" />
                    <SPLIT distance="150" swimtime="00:01:42.52" />
                    <SPLIT distance="175" swimtime="00:02:00.59" />
                    <SPLIT distance="200" swimtime="00:02:18.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106981" lastname="STEENBERGEN" firstname="Marrit" gender="F" birthdate="2000-01-11">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:51.92" eventid="13" heat="9" lane="3">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.75" eventid="43" heat="4" lane="5">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.15" eventid="6" heat="5" lane="6">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:00:58.15" eventid="22" heat="2" lane="4">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="3" lane="6" heat="1" heatid="10113" swimtime="00:00:51.25" reactiontime="+73" points="942">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.77" />
                    <SPLIT distance="50" swimtime="00:00:24.66" />
                    <SPLIT distance="75" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:00:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="2" lane="3" heat="9" heatid="90013" swimtime="00:00:52.23" reactiontime="+75" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.01" />
                    <SPLIT distance="50" swimtime="00:00:25.19" />
                    <SPLIT distance="75" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="4" lane="4" heat="1" heatid="10213" swimtime="00:00:51.85" reactiontime="+73" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                    <SPLIT distance="75" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:00:51.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="143" place="3" lane="4" heat="1" heatid="10143" swimtime="00:01:52.28" reactiontime="+73" points="948">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.25" />
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                    <SPLIT distance="75" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:00:54.59" />
                    <SPLIT distance="125" swimtime="00:01:08.83" />
                    <SPLIT distance="150" swimtime="00:01:23.42" />
                    <SPLIT distance="175" swimtime="00:01:38.05" />
                    <SPLIT distance="200" swimtime="00:01:52.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="1" lane="5" heat="4" heatid="40043" swimtime="00:01:52.83" reactiontime="+72" points="934">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.14" />
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="75" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:00:54.03" />
                    <SPLIT distance="125" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:23.05" />
                    <SPLIT distance="175" swimtime="00:01:38.13" />
                    <SPLIT distance="200" swimtime="00:01:52.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106" place="4" lane="3" heat="1" heatid="10106" swimtime="00:02:04.94" reactiontime="+73" points="927">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                    <SPLIT distance="75" swimtime="00:00:43.07" />
                    <SPLIT distance="100" swimtime="00:00:58.56" />
                    <SPLIT distance="125" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:35.32" />
                    <SPLIT distance="175" swimtime="00:01:50.79" />
                    <SPLIT distance="200" swimtime="00:02:04.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="3" lane="6" heat="5" heatid="50006" swimtime="00:02:06.01" reactiontime="+73" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:27.13" />
                    <SPLIT distance="75" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:00:59.56" />
                    <SPLIT distance="125" swimtime="00:01:17.37" />
                    <SPLIT distance="150" swimtime="00:01:36.00" />
                    <SPLIT distance="175" swimtime="00:01:51.40" />
                    <SPLIT distance="200" swimtime="00:02:06.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="1" lane="4" heat="1" heatid="10122" swimtime="00:00:57.53" reactiontime="+57" points="947">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                    <SPLIT distance="75" swimtime="00:00:43.53" />
                    <SPLIT distance="100" swimtime="00:00:57.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="2" lane="4" heat="2" heatid="20022" swimtime="00:00:58.87" reactiontime="+74" points="884">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="75" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:00:58.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="1" lane="4" heat="1" heatid="10222" swimtime="00:00:57.65" reactiontime="+73" points="941">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:26.52" />
                    <SPLIT distance="75" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:00:57.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109023" lastname="BUSCH" firstname="Kim" gender="F" birthdate="1998-06-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.17" eventid="13" heat="8" lane="7">
                  <MEETINFO date="2021-09-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:24.15" eventid="30" heat="7" lane="2">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="23" lane="7" heat="8" heatid="80013" swimtime="00:00:53.84" reactiontime="+76" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                    <SPLIT distance="75" swimtime="00:00:39.40" />
                    <SPLIT distance="100" swimtime="00:00:53.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="14" lane="2" heat="7" heatid="70030" swimtime="00:00:24.37" reactiontime="+72" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="14" lane="1" heat="1" heatid="10230" swimtime="00:00:24.34" reactiontime="+75" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:24.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109036" lastname="VERMEULEN" firstname="Tessa" gender="F" birthdate="1998-01-29">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.34" eventid="45" heat="5" lane="7">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="20" lane="7" heat="5" heatid="50045" swimtime="00:02:06.58" reactiontime="+63" points="829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="75" swimtime="00:00:45.35" />
                    <SPLIT distance="100" swimtime="00:01:01.37" />
                    <SPLIT distance="125" swimtime="00:01:17.32" />
                    <SPLIT distance="150" swimtime="00:01:33.81" />
                    <SPLIT distance="175" swimtime="00:01:50.26" />
                    <SPLIT distance="200" swimtime="00:02:06.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154332" lastname="DE JONG" firstname="Imani" gender="F" birthdate="2002-05-28">
              <ENTRIES>
                <ENTRY entrytime="00:04:05.68" eventid="1" heat="4" lane="8">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:08:28.90" eventid="12" heat="2" lane="6">
                  <MEETINFO date="2021-10-03" />
                </ENTRY>
                <ENTRY entrytime="00:16:19.04" eventid="33" heat="2" lane="3">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="11" lane="8" heat="4" heatid="40001" swimtime="00:04:04.65" reactiontime="+71" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.93" />
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                    <SPLIT distance="75" swimtime="00:00:42.94" />
                    <SPLIT distance="100" swimtime="00:00:58.35" />
                    <SPLIT distance="125" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:01:29.15" />
                    <SPLIT distance="175" swimtime="00:01:44.70" />
                    <SPLIT distance="200" swimtime="00:02:00.07" />
                    <SPLIT distance="225" swimtime="00:02:15.65" />
                    <SPLIT distance="250" swimtime="00:02:31.31" />
                    <SPLIT distance="275" swimtime="00:02:47.05" />
                    <SPLIT distance="300" swimtime="00:03:02.68" />
                    <SPLIT distance="325" swimtime="00:03:18.48" />
                    <SPLIT distance="350" swimtime="00:03:34.26" />
                    <SPLIT distance="375" swimtime="00:03:49.65" />
                    <SPLIT distance="400" swimtime="00:04:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="10" lane="6" heat="2" heatid="20012" swimtime="00:08:25.84" reactiontime="+71" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                    <SPLIT distance="75" swimtime="00:00:44.01" />
                    <SPLIT distance="100" swimtime="00:00:59.80" />
                    <SPLIT distance="125" swimtime="00:01:15.53" />
                    <SPLIT distance="150" swimtime="00:01:31.38" />
                    <SPLIT distance="175" swimtime="00:01:47.25" />
                    <SPLIT distance="200" swimtime="00:02:03.14" />
                    <SPLIT distance="225" swimtime="00:02:19.05" />
                    <SPLIT distance="250" swimtime="00:02:34.94" />
                    <SPLIT distance="275" swimtime="00:02:51.01" />
                    <SPLIT distance="300" swimtime="00:03:07.02" />
                    <SPLIT distance="325" swimtime="00:03:23.04" />
                    <SPLIT distance="350" swimtime="00:03:39.14" />
                    <SPLIT distance="375" swimtime="00:03:55.19" />
                    <SPLIT distance="400" swimtime="00:04:11.17" />
                    <SPLIT distance="425" swimtime="00:04:27.17" />
                    <SPLIT distance="450" swimtime="00:04:43.29" />
                    <SPLIT distance="475" swimtime="00:04:59.31" />
                    <SPLIT distance="500" swimtime="00:05:15.42" />
                    <SPLIT distance="525" swimtime="00:05:31.47" />
                    <SPLIT distance="550" swimtime="00:05:47.64" />
                    <SPLIT distance="575" swimtime="00:06:03.78" />
                    <SPLIT distance="600" swimtime="00:06:19.77" />
                    <SPLIT distance="625" swimtime="00:06:35.68" />
                    <SPLIT distance="650" swimtime="00:06:51.65" />
                    <SPLIT distance="675" swimtime="00:07:07.58" />
                    <SPLIT distance="700" swimtime="00:07:23.63" />
                    <SPLIT distance="725" swimtime="00:07:39.71" />
                    <SPLIT distance="750" swimtime="00:07:55.71" />
                    <SPLIT distance="775" swimtime="00:08:11.13" />
                    <SPLIT distance="800" swimtime="00:08:25.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="10" lane="3" heat="2" heatid="20033" swimtime="00:16:15.61" reactiontime="+73" points="833">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:28.52" />
                    <SPLIT distance="75" swimtime="00:00:44.06" />
                    <SPLIT distance="100" swimtime="00:01:00.00" />
                    <SPLIT distance="125" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:31.95" />
                    <SPLIT distance="175" swimtime="00:01:47.89" />
                    <SPLIT distance="200" swimtime="00:02:04.05" />
                    <SPLIT distance="225" swimtime="00:02:20.10" />
                    <SPLIT distance="250" swimtime="00:02:36.11" />
                    <SPLIT distance="275" swimtime="00:02:52.35" />
                    <SPLIT distance="300" swimtime="00:03:08.53" />
                    <SPLIT distance="325" swimtime="00:03:24.61" />
                    <SPLIT distance="350" swimtime="00:03:40.76" />
                    <SPLIT distance="375" swimtime="00:03:56.91" />
                    <SPLIT distance="400" swimtime="00:04:13.02" />
                    <SPLIT distance="425" swimtime="00:04:29.15" />
                    <SPLIT distance="450" swimtime="00:04:45.38" />
                    <SPLIT distance="475" swimtime="00:05:01.60" />
                    <SPLIT distance="500" swimtime="00:05:17.79" />
                    <SPLIT distance="525" swimtime="00:05:34.01" />
                    <SPLIT distance="550" swimtime="00:05:50.25" />
                    <SPLIT distance="575" swimtime="00:06:06.60" />
                    <SPLIT distance="600" swimtime="00:06:22.92" />
                    <SPLIT distance="625" swimtime="00:06:39.31" />
                    <SPLIT distance="650" swimtime="00:06:55.60" />
                    <SPLIT distance="675" swimtime="00:07:11.98" />
                    <SPLIT distance="700" swimtime="00:07:28.40" />
                    <SPLIT distance="725" swimtime="00:07:44.81" />
                    <SPLIT distance="750" swimtime="00:08:01.25" />
                    <SPLIT distance="775" swimtime="00:08:17.83" />
                    <SPLIT distance="800" swimtime="00:08:34.15" />
                    <SPLIT distance="825" swimtime="00:08:50.74" />
                    <SPLIT distance="850" swimtime="00:09:07.16" />
                    <SPLIT distance="875" swimtime="00:09:23.92" />
                    <SPLIT distance="900" swimtime="00:09:40.42" />
                    <SPLIT distance="925" swimtime="00:09:57.09" />
                    <SPLIT distance="950" swimtime="00:10:13.63" />
                    <SPLIT distance="975" swimtime="00:10:30.10" />
                    <SPLIT distance="1000" swimtime="00:10:46.59" />
                    <SPLIT distance="1025" swimtime="00:11:03.21" />
                    <SPLIT distance="1050" swimtime="00:11:19.77" />
                    <SPLIT distance="1075" swimtime="00:11:36.40" />
                    <SPLIT distance="1100" swimtime="00:11:52.92" />
                    <SPLIT distance="1125" swimtime="00:12:09.39" />
                    <SPLIT distance="1150" swimtime="00:12:25.83" />
                    <SPLIT distance="1175" swimtime="00:12:42.31" />
                    <SPLIT distance="1200" swimtime="00:12:58.70" />
                    <SPLIT distance="1225" swimtime="00:13:15.06" />
                    <SPLIT distance="1250" swimtime="00:13:31.48" />
                    <SPLIT distance="1275" swimtime="00:13:47.73" />
                    <SPLIT distance="1300" swimtime="00:14:04.06" />
                    <SPLIT distance="1325" swimtime="00:14:20.43" />
                    <SPLIT distance="1350" swimtime="00:14:36.90" />
                    <SPLIT distance="1375" swimtime="00:14:53.39" />
                    <SPLIT distance="1400" swimtime="00:15:09.96" />
                    <SPLIT distance="1425" swimtime="00:15:26.52" />
                    <SPLIT distance="1450" swimtime="00:15:43.15" />
                    <SPLIT distance="1475" swimtime="00:15:59.55" />
                    <SPLIT distance="1500" swimtime="00:16:15.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154337" lastname="HOLKENBORG" firstname="Silke" gender="F" birthdate="2001-08-31">
              <ENTRIES>
                <ENTRY entrytime="00:04:06.79" eventid="1" heat="3" lane="8">
                  <MEETINFO date="2022-07-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="16" lane="8" heat="3" heatid="30001" swimtime="00:04:08.75" reactiontime="+68" points="831">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="75" swimtime="00:00:44.07" />
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="125" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:01:31.06" />
                    <SPLIT distance="175" swimtime="00:01:46.96" />
                    <SPLIT distance="200" swimtime="00:02:02.83" />
                    <SPLIT distance="225" swimtime="00:02:18.66" />
                    <SPLIT distance="250" swimtime="00:02:34.43" />
                    <SPLIT distance="275" swimtime="00:02:50.42" />
                    <SPLIT distance="300" swimtime="00:03:06.33" />
                    <SPLIT distance="325" swimtime="00:03:22.08" />
                    <SPLIT distance="350" swimtime="00:03:37.72" />
                    <SPLIT distance="375" swimtime="00:03:53.57" />
                    <SPLIT distance="400" swimtime="00:04:08.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130232" lastname="VAN ROON" firstname="Valerie" gender="F" birthdate="1998-08-13">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:23.94" eventid="30" heat="6" lane="3">
                  <MEETINFO date="2022-07-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="30" place="12" lane="3" heat="6" heatid="60030" swimtime="00:00:24.33" reactiontime="+67" points="837">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.77" />
                    <SPLIT distance="50" swimtime="00:00:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="10" lane="7" heat="1" heatid="10230" swimtime="00:00:24.19" reactiontime="+69" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:24.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Netherlands">
              <RESULTS>
                <RESULT eventid="109" place="8" lane="7" heat="1" swimtime="00:03:08.84" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.56" />
                    <SPLIT distance="50" swimtime="00:00:22.75" />
                    <SPLIT distance="75" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:00:47.74" />
                    <SPLIT distance="125" swimtime="00:00:57.84" />
                    <SPLIT distance="150" swimtime="00:01:09.68" />
                    <SPLIT distance="175" swimtime="00:01:22.03" />
                    <SPLIT distance="200" swimtime="00:01:34.49" />
                    <SPLIT distance="225" swimtime="00:01:44.26" />
                    <SPLIT distance="250" swimtime="00:01:56.26" />
                    <SPLIT distance="275" swimtime="00:02:08.59" />
                    <SPLIT distance="300" swimtime="00:02:21.45" />
                    <SPLIT distance="325" swimtime="00:02:31.32" />
                    <SPLIT distance="350" swimtime="00:02:43.21" />
                    <SPLIT distance="375" swimtime="00:02:55.84" />
                    <SPLIT distance="400" swimtime="00:03:08.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109044" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="154353" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="106982" reactiontime="+13" />
                    <RELAYPOSITION number="4" athleteid="129673" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="6" lane="5" heat="2" swimtime="00:03:08.58" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.47" />
                    <SPLIT distance="50" swimtime="00:00:22.48" />
                    <SPLIT distance="75" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:00:47.24" />
                    <SPLIT distance="125" swimtime="00:00:57.36" />
                    <SPLIT distance="150" swimtime="00:01:09.26" />
                    <SPLIT distance="175" swimtime="00:01:21.79" />
                    <SPLIT distance="200" swimtime="00:01:34.55" />
                    <SPLIT distance="225" swimtime="00:01:44.73" />
                    <SPLIT distance="250" swimtime="00:01:56.57" />
                    <SPLIT distance="275" swimtime="00:02:08.78" />
                    <SPLIT distance="300" swimtime="00:02:21.07" />
                    <SPLIT distance="325" swimtime="00:02:31.61" />
                    <SPLIT distance="350" swimtime="00:02:43.50" />
                    <SPLIT distance="375" swimtime="00:02:56.09" />
                    <SPLIT distance="400" swimtime="00:03:08.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109044" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="154357" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="154353" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="154356" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Netherlands">
              <RESULTS>
                <RESULT eventid="48" place="11" lane="3" heat="3" swimtime="00:03:28.61" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                    <SPLIT distance="50" swimtime="00:00:25.77" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:54.41" />
                    <SPLIT distance="125" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:20.83" />
                    <SPLIT distance="175" swimtime="00:01:36.23" />
                    <SPLIT distance="200" swimtime="00:01:51.75" />
                    <SPLIT distance="225" swimtime="00:02:02.01" />
                    <SPLIT distance="250" swimtime="00:02:14.74" />
                    <SPLIT distance="275" swimtime="00:02:28.17" />
                    <SPLIT distance="300" swimtime="00:02:41.87" />
                    <SPLIT distance="325" swimtime="00:02:51.79" />
                    <SPLIT distance="350" swimtime="00:03:03.55" />
                    <SPLIT distance="375" swimtime="00:03:16.01" />
                    <SPLIT distance="400" swimtime="00:03:28.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109044" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="154353" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="106982" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="154357" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Netherlands">
              <RESULTS>
                <RESULT eventid="126" place="3" lane="4" heat="1" swimtime="00:01:23.75" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.09" />
                    <SPLIT distance="50" swimtime="00:00:21.24" />
                    <SPLIT distance="75" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:00:42.08" />
                    <SPLIT distance="125" swimtime="00:00:51.81" />
                    <SPLIT distance="150" swimtime="00:01:03.03" />
                    <SPLIT distance="175" swimtime="00:01:12.66" />
                    <SPLIT distance="200" swimtime="00:01:23.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154357" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="106982" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="109044" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="129673" reactiontime="+4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="1" lane="4" heat="2" swimtime="00:01:23.70" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:21.28" />
                    <SPLIT distance="75" swimtime="00:00:30.88" />
                    <SPLIT distance="100" swimtime="00:00:42.07" />
                    <SPLIT distance="125" swimtime="00:00:51.89" />
                    <SPLIT distance="150" swimtime="00:01:03.14" />
                    <SPLIT distance="175" swimtime="00:01:12.62" />
                    <SPLIT distance="200" swimtime="00:01:23.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154357" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="106982" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="109044" reactiontime="+22" />
                    <RELAYPOSITION number="4" athleteid="129673" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Netherlands">
              <RESULTS>
                <RESULT eventid="127" place="3" lane="3" heat="1" swimtime="00:01:28.53" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.05" />
                    <SPLIT distance="50" swimtime="00:00:21.14" />
                    <SPLIT distance="75" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:00:41.75" />
                    <SPLIT distance="125" swimtime="00:00:52.73" />
                    <SPLIT distance="150" swimtime="00:01:05.10" />
                    <SPLIT distance="175" swimtime="00:01:16.37" />
                    <SPLIT distance="200" swimtime="00:01:28.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154357" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="129673" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="109026" reactiontime="+10" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="3" lane="4" heat="3" swimtime="00:01:29.95" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.44" />
                    <SPLIT distance="50" swimtime="00:00:21.71" />
                    <SPLIT distance="75" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:00:42.67" />
                    <SPLIT distance="125" swimtime="00:00:53.77" />
                    <SPLIT distance="150" swimtime="00:01:06.28" />
                    <SPLIT distance="175" swimtime="00:01:17.62" />
                    <SPLIT distance="200" swimtime="00:01:29.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109044" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="106982" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="109026" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Netherlands">
              <RESULTS>
                <RESULT eventid="108" place="5" lane="5" heat="1" swimtime="00:03:29.59" reactiontime="+75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                    <SPLIT distance="75" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:00:53.37" />
                    <SPLIT distance="125" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:18.33" />
                    <SPLIT distance="175" swimtime="00:01:31.85" />
                    <SPLIT distance="200" swimtime="00:01:45.70" />
                    <SPLIT distance="225" swimtime="00:01:57.32" />
                    <SPLIT distance="250" swimtime="00:02:10.58" />
                    <SPLIT distance="275" swimtime="00:02:24.62" />
                    <SPLIT distance="300" swimtime="00:02:38.68" />
                    <SPLIT distance="325" swimtime="00:02:50.18" />
                    <SPLIT distance="350" swimtime="00:03:03.32" />
                    <SPLIT distance="375" swimtime="00:03:16.41" />
                    <SPLIT distance="400" swimtime="00:03:29.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109023" reactiontime="+75" />
                    <RELAYPOSITION number="2" athleteid="109025" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="130232" reactiontime="+43" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="2" lane="5" heat="1" swimtime="00:03:30.42" reactiontime="+73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.95" />
                    <SPLIT distance="50" swimtime="00:00:25.06" />
                    <SPLIT distance="75" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:00:53.28" />
                    <SPLIT distance="125" swimtime="00:01:04.90" />
                    <SPLIT distance="150" swimtime="00:01:18.12" />
                    <SPLIT distance="175" swimtime="00:01:32.08" />
                    <SPLIT distance="200" swimtime="00:01:46.40" />
                    <SPLIT distance="225" swimtime="00:01:58.06" />
                    <SPLIT distance="250" swimtime="00:02:11.35" />
                    <SPLIT distance="275" swimtime="00:02:24.96" />
                    <SPLIT distance="300" swimtime="00:02:38.70" />
                    <SPLIT distance="325" swimtime="00:02:50.36" />
                    <SPLIT distance="350" swimtime="00:03:03.51" />
                    <SPLIT distance="375" swimtime="00:03:17.05" />
                    <SPLIT distance="400" swimtime="00:03:30.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109023" reactiontime="+73" />
                    <RELAYPOSITION number="2" athleteid="130232" reactiontime="+35" />
                    <RELAYPOSITION number="3" athleteid="109025" reactiontime="+21" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Netherlands">
              <RESULTS>
                <RESULT eventid="147" place="4" lane="7" heat="1" swimtime="00:03:47.70" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="75" swimtime="00:00:41.93" />
                    <SPLIT distance="100" swimtime="00:00:56.53" />
                    <SPLIT distance="125" swimtime="00:01:10.37" />
                    <SPLIT distance="150" swimtime="00:01:26.97" />
                    <SPLIT distance="175" swimtime="00:01:44.27" />
                    <SPLIT distance="200" swimtime="00:02:01.81" />
                    <SPLIT distance="225" swimtime="00:02:13.02" />
                    <SPLIT distance="250" swimtime="00:02:27.13" />
                    <SPLIT distance="275" swimtime="00:02:41.82" />
                    <SPLIT distance="300" swimtime="00:02:57.23" />
                    <SPLIT distance="325" swimtime="00:03:08.47" />
                    <SPLIT distance="350" swimtime="00:03:21.51" />
                    <SPLIT distance="375" swimtime="00:03:34.70" />
                    <SPLIT distance="400" swimtime="00:03:47.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109025" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="129677" reactiontime="+27" />
                    <RELAYPOSITION number="3" athleteid="109026" reactiontime="+15" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+11" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="6" lane="6" heat="2" swimtime="00:03:52.95" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="75" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:00:56.78" />
                    <SPLIT distance="125" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:27.00" />
                    <SPLIT distance="175" swimtime="00:01:44.03" />
                    <SPLIT distance="200" swimtime="00:02:01.53" />
                    <SPLIT distance="225" swimtime="00:02:13.14" />
                    <SPLIT distance="250" swimtime="00:02:27.22" />
                    <SPLIT distance="275" swimtime="00:02:42.40" />
                    <SPLIT distance="300" swimtime="00:02:59.34" />
                    <SPLIT distance="325" swimtime="00:03:11.38" />
                    <SPLIT distance="350" swimtime="00:03:24.73" />
                    <SPLIT distance="375" swimtime="00:03:38.85" />
                    <SPLIT distance="400" swimtime="00:03:52.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109026" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="129677" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="109023" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="130232" reactiontime="+58" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Netherlands">
              <RESULTS>
                <RESULT eventid="117" place="4" lane="3" heat="1" swimtime="00:07:40.54" reactiontime="+73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.79" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="75" swimtime="00:00:41.35" />
                    <SPLIT distance="100" swimtime="00:00:55.99" />
                    <SPLIT distance="125" swimtime="00:01:10.90" />
                    <SPLIT distance="150" swimtime="00:01:26.23" />
                    <SPLIT distance="175" swimtime="00:01:41.63" />
                    <SPLIT distance="200" swimtime="00:01:56.88" />
                    <SPLIT distance="225" swimtime="00:02:08.66" />
                    <SPLIT distance="250" swimtime="00:02:22.13" />
                    <SPLIT distance="275" swimtime="00:02:36.29" />
                    <SPLIT distance="300" swimtime="00:02:50.58" />
                    <SPLIT distance="325" swimtime="00:03:04.81" />
                    <SPLIT distance="350" swimtime="00:03:19.49" />
                    <SPLIT distance="375" swimtime="00:03:34.18" />
                    <SPLIT distance="400" swimtime="00:03:48.82" />
                    <SPLIT distance="425" swimtime="00:04:01.17" />
                    <SPLIT distance="450" swimtime="00:04:15.36" />
                    <SPLIT distance="475" swimtime="00:04:30.01" />
                    <SPLIT distance="500" swimtime="00:04:44.95" />
                    <SPLIT distance="525" swimtime="00:04:59.94" />
                    <SPLIT distance="550" swimtime="00:05:15.05" />
                    <SPLIT distance="575" swimtime="00:05:30.21" />
                    <SPLIT distance="600" swimtime="00:05:44.90" />
                    <SPLIT distance="625" swimtime="00:05:56.89" />
                    <SPLIT distance="650" swimtime="00:06:10.85" />
                    <SPLIT distance="675" swimtime="00:06:25.55" />
                    <SPLIT distance="700" swimtime="00:06:40.31" />
                    <SPLIT distance="725" swimtime="00:06:55.27" />
                    <SPLIT distance="750" swimtime="00:07:10.37" />
                    <SPLIT distance="775" swimtime="00:07:25.62" />
                    <SPLIT distance="800" swimtime="00:07:40.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109036" reactiontime="+73" />
                    <RELAYPOSITION number="2" athleteid="106981" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="154337" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="154332" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="3" lane="3" heat="1" swimtime="00:07:45.73" reactiontime="+73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:26.86" />
                    <SPLIT distance="75" swimtime="00:00:41.27" />
                    <SPLIT distance="100" swimtime="00:00:55.95" />
                    <SPLIT distance="125" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:25.81" />
                    <SPLIT distance="175" swimtime="00:01:41.44" />
                    <SPLIT distance="200" swimtime="00:01:56.89" />
                    <SPLIT distance="225" swimtime="00:02:09.36" />
                    <SPLIT distance="250" swimtime="00:02:23.50" />
                    <SPLIT distance="275" swimtime="00:02:38.40" />
                    <SPLIT distance="300" swimtime="00:02:53.57" />
                    <SPLIT distance="325" swimtime="00:03:09.02" />
                    <SPLIT distance="350" swimtime="00:03:24.47" />
                    <SPLIT distance="375" swimtime="00:03:39.99" />
                    <SPLIT distance="400" swimtime="00:03:54.94" />
                    <SPLIT distance="425" swimtime="00:04:07.61" />
                    <SPLIT distance="450" swimtime="00:04:21.80" />
                    <SPLIT distance="475" swimtime="00:04:36.18" />
                    <SPLIT distance="500" swimtime="00:04:50.99" />
                    <SPLIT distance="525" swimtime="00:05:05.81" />
                    <SPLIT distance="550" swimtime="00:05:20.61" />
                    <SPLIT distance="575" swimtime="00:05:35.87" />
                    <SPLIT distance="600" swimtime="00:05:50.57" />
                    <SPLIT distance="625" swimtime="00:06:02.48" />
                    <SPLIT distance="650" swimtime="00:06:16.52" />
                    <SPLIT distance="675" swimtime="00:06:31.08" />
                    <SPLIT distance="700" swimtime="00:06:46.03" />
                    <SPLIT distance="725" swimtime="00:07:01.05" />
                    <SPLIT distance="750" swimtime="00:07:16.31" />
                    <SPLIT distance="775" swimtime="00:07:31.24" />
                    <SPLIT distance="800" swimtime="00:07:45.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109036" reactiontime="+73" />
                    <RELAYPOSITION number="2" athleteid="154332" reactiontime="+60" />
                    <RELAYPOSITION number="3" athleteid="154337" reactiontime="+48" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+36" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Netherlands">
              <RESULTS>
                <RESULT eventid="125" place="3" lane="6" heat="1" swimtime="00:01:35.36" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:24.20" />
                    <SPLIT distance="75" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:00:47.67" />
                    <SPLIT distance="125" swimtime="00:00:59.00" />
                    <SPLIT distance="150" swimtime="00:01:11.68" />
                    <SPLIT distance="175" swimtime="00:01:22.90" />
                    <SPLIT distance="200" swimtime="00:01:35.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109023" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="109026" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="109025" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="130232" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="4" lane="5" heat="2" swimtime="00:01:36.32" reactiontime="+77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:24.06" />
                    <SPLIT distance="75" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:00:47.71" />
                    <SPLIT distance="125" swimtime="00:00:59.00" />
                    <SPLIT distance="150" swimtime="00:01:11.46" />
                    <SPLIT distance="175" swimtime="00:01:23.38" />
                    <SPLIT distance="200" swimtime="00:01:36.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109023" reactiontime="+77" />
                    <RELAYPOSITION number="2" athleteid="109026" reactiontime="+30" />
                    <RELAYPOSITION number="3" athleteid="130232" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="109036" reactiontime="+34" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Netherlands">
              <RESULTS>
                <RESULT eventid="134" place="5" lane="2" heat="1" swimtime="00:01:43.72" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                    <SPLIT distance="75" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:00:56.01" />
                    <SPLIT distance="125" swimtime="00:01:06.97" />
                    <SPLIT distance="150" swimtime="00:01:20.40" />
                    <SPLIT distance="175" swimtime="00:01:31.51" />
                    <SPLIT distance="200" swimtime="00:01:43.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109025" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="129677" reactiontime="+11" />
                    <RELAYPOSITION number="3" athleteid="109026" reactiontime="+17" />
                    <RELAYPOSITION number="4" athleteid="106981" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="5" lane="5" heat="2" swimtime="00:01:46.06" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                    <SPLIT distance="75" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:00:56.45" />
                    <SPLIT distance="125" swimtime="00:01:08.13" />
                    <SPLIT distance="150" swimtime="00:01:21.86" />
                    <SPLIT distance="175" swimtime="00:01:33.47" />
                    <SPLIT distance="200" swimtime="00:01:46.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109025" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="129677" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="109023" reactiontime="+58" />
                    <RELAYPOSITION number="4" athleteid="130232" reactiontime="+44" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Netherlands">
              <RESULTS>
                <RESULT eventid="111" place="-1" lane="6" heat="1" status="DSQ" swimtime="00:01:36.40" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                    <SPLIT distance="75" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:00:51.56" />
                    <SPLIT distance="125" swimtime="00:01:02.60" />
                    <SPLIT distance="150" swimtime="00:01:16.06" />
                    <SPLIT distance="175" swimtime="00:01:25.39" />
                    <SPLIT distance="200" swimtime="00:01:36.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109025" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="154353" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="109026" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="129673" reactiontime="-4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="4" lane="4" heat="4" swimtime="00:01:38.59" reactiontime="+51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:26.37" />
                    <SPLIT distance="75" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:00:52.63" />
                    <SPLIT distance="125" swimtime="00:01:02.56" />
                    <SPLIT distance="150" swimtime="00:01:14.76" />
                    <SPLIT distance="175" swimtime="00:01:26.09" />
                    <SPLIT distance="200" swimtime="00:01:38.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109025" reactiontime="+51" />
                    <RELAYPOSITION number="2" athleteid="154353" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="106982" reactiontime="+30" />
                    <RELAYPOSITION number="4" athleteid="130232" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Netherlands">
              <RESULTS>
                <RESULT eventid="135" place="8" lane="7" heat="1" swimtime="00:01:33.43" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.05" />
                    <SPLIT distance="75" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:00:50.32" />
                    <SPLIT distance="125" swimtime="00:01:00.18" />
                    <SPLIT distance="150" swimtime="00:01:12.59" />
                    <SPLIT distance="175" swimtime="00:01:22.18" />
                    <SPLIT distance="200" swimtime="00:01:33.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109044" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="154353" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="106982" reactiontime="+21" />
                    <RELAYPOSITION number="4" athleteid="129673" reactiontime="+3" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="6" lane="2" heat="1" swimtime="00:01:33.20" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.60" />
                    <SPLIT distance="50" swimtime="00:00:23.89" />
                    <SPLIT distance="75" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:00:49.97" />
                    <SPLIT distance="125" swimtime="00:00:59.83" />
                    <SPLIT distance="150" swimtime="00:01:12.25" />
                    <SPLIT distance="175" swimtime="00:01:21.98" />
                    <SPLIT distance="200" swimtime="00:01:33.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="109044" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="154353" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="106982" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="154357" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Nepal" shortname="NEP" code="NEP" nation="NEP" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="183417" lastname="KUMAL" firstname="Bikash" gender="M" birthdate="2004-04-25">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.94" eventid="16" heat="1" lane="5">
                  <MEETINFO date="2022-08-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.50" eventid="41" heat="2" lane="3">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="57" lane="5" heat="1" heatid="10016" swimtime="00:01:07.50" reactiontime="+62" points="549">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.61" />
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="75" swimtime="00:00:49.52" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="54" lane="3" heat="2" heatid="20041" swimtime="00:00:31.11" reactiontime="+64" points="515">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.28" />
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214408" lastname="SHRESTHA" firstname="Ervin" gender="M" birthdate="2007-08-05">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="14" heat="1" lane="2" />
                <ENTRY entrytime="NT" eventid="44" heat="1" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="79" lane="2" heat="1" heatid="10014" swimtime="00:00:56.87" reactiontime="+71" points="490">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.32" />
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                    <SPLIT distance="75" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:00:56.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="46" lane="1" heat="1" heatid="10044" swimtime="00:02:05.03" reactiontime="+70" points="502">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                    <SPLIT distance="75" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:01:00.22" />
                    <SPLIT distance="125" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:01:32.72" />
                    <SPLIT distance="175" swimtime="00:01:49.25" />
                    <SPLIT distance="200" swimtime="00:02:05.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197746" lastname="TANDUKAR" firstname="Anushiya" gender="F" birthdate="2006-03-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.77" eventid="13" heat="3" lane="1">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.03" eventid="30" heat="2" lane="4">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="56" lane="1" heat="3" heatid="30013" swimtime="00:01:02.49" reactiontime="+77" points="519">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="75" swimtime="00:00:46.60" />
                    <SPLIT distance="100" swimtime="00:01:02.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="47" lane="4" heat="2" heatid="20030" swimtime="00:00:28.92" reactiontime="+70" points="498">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214407" lastname="NEUPANE" firstname="Rosha" gender="F" birthdate="2007-08-05">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="18" heat="1" lane="5" />
                <ENTRY entrytime="NT" eventid="4" heat="1" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="49" lane="5" heat="1" heatid="10018" swimtime="00:00:35.28" reactiontime="+81" points="367">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.62" />
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="39" lane="6" heat="1" heatid="10004" swimtime="00:00:31.95" reactiontime="+79" points="444">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.68" />
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Nigeria" shortname="NGR" code="NGR" nation="NGR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="196654" lastname="OPUTE" firstname="Clinton" gender="M" birthdate="2003-04-11">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.02" eventid="14" heat="1" lane="4">
                  <MEETINFO date="2021-10-14" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.14" eventid="31" heat="4" lane="8">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="73" lane="4" heat="1" heatid="10014" swimtime="00:00:53.66" reactiontime="+66" points="583">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:25.39" />
                    <SPLIT distance="75" swimtime="00:00:39.36" />
                    <SPLIT distance="100" swimtime="00:00:53.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="62" lane="8" heat="4" heatid="40031" swimtime="00:00:24.47" reactiontime="+68" points="559">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:24.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Niger" shortname="NIG" code="NIG" nation="NIG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="122970" lastname="SEYDOU LANCINA" firstname="Alassane" gender="M" birthdate="1993-09-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.28" eventid="5" heat="3" lane="6">
                  <MEETINFO date="2022-08-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.61" eventid="31" heat="5" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="57" lane="6" heat="3" heatid="30005" swimtime="00:00:26.63" reactiontime="+81" points="544">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:26.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="53" lane="1" heat="5" heatid="50031" swimtime="00:00:23.64" reactiontime="+75" points="620">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.67" />
                    <SPLIT distance="50" swimtime="00:00:23.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154815" lastname="AHMADOU YOUSSOUFOU" firstname="Salima" gender="F" birthdate="2003-10-21">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="15" heat="1" lane="3" />
                <ENTRY entrytime="00:00:55.67" eventid="40" heat="2" lane="7">
                  <MEETINFO date="2021-10-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="52" lane="3" heat="1" heatid="10015" swimtime="00:01:58.58" reactiontime="+76" points="145">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.33" />
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                    <SPLIT distance="75" swimtime="00:01:23.11" />
                    <SPLIT distance="100" swimtime="00:01:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="44" lane="7" heat="2" heatid="20040" swimtime="00:00:48.33" reactiontime="+66" points="206">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.46" />
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Northern Mariana Islands" shortname="NMA" code="NMA" nation="NMA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="214457" lastname="ALEKSENKO" firstname="Isaiah" gender="M" birthdate="2006-05-06">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="39" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="21" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="41" lane="4" heat="1" heatid="10039" swimtime="00:00:54.55" reactiontime="+61" points="671">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:25.29" />
                    <SPLIT distance="75" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:00:54.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="24" lane="3" heat="1" heatid="10021" swimtime="00:02:02.96" reactiontime="+63" points="682">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                    <SPLIT distance="75" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:00:56.65" />
                    <SPLIT distance="125" swimtime="00:01:12.61" />
                    <SPLIT distance="150" swimtime="00:01:29.06" />
                    <SPLIT distance="175" swimtime="00:01:46.01" />
                    <SPLIT distance="200" swimtime="00:02:02.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161275" lastname="SUZUKI" firstname="Jinnosuke" gender="M" birthdate="2005-10-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.72" eventid="14" heat="3" lane="6">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.27" eventid="44" heat="1" lane="3">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="75" lane="6" heat="3" heatid="30014" swimtime="00:00:54.48" reactiontime="+62" points="557">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.48" />
                    <SPLIT distance="50" swimtime="00:00:25.95" />
                    <SPLIT distance="75" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:00:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="43" lane="3" heat="1" heatid="10044" swimtime="00:01:56.27" reactiontime="+63" points="624">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                    <SPLIT distance="75" swimtime="00:00:41.23" />
                    <SPLIT distance="100" swimtime="00:00:55.92" />
                    <SPLIT distance="125" swimtime="00:01:10.68" />
                    <SPLIT distance="150" swimtime="00:01:25.82" />
                    <SPLIT distance="175" swimtime="00:01:41.04" />
                    <SPLIT distance="200" swimtime="00:01:56.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197310" lastname="LITULUMAR" firstname="Shoko" gender="F" birthdate="2007-01-27">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="2" heat="1" lane="8" />
                <ENTRY entrytime="00:00:33.85" eventid="18" heat="2" lane="3">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="46" lane="8" heat="1" heatid="10002" swimtime="00:01:14.72" reactiontime="+63" points="396">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:35.63" />
                    <SPLIT distance="75" swimtime="00:00:55.21" />
                    <SPLIT distance="100" swimtime="00:01:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="46" lane="3" heat="2" heatid="20018" swimtime="00:00:33.86" reactiontime="+60" points="415">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.62" />
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201852" lastname="BATALLONES" firstname="Maria Corazon Ayson" gender="F" birthdate="2008-06-03">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:26.01" eventid="15" heat="1" lane="4">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:37.77" eventid="40" heat="2" lane="4">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="49" lane="4" heat="1" heatid="10015" swimtime="00:01:18.08" reactiontime="+63" points="509">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.07" />
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="75" swimtime="00:00:57.26" />
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="36" lane="4" heat="2" heatid="20040" swimtime="00:00:34.58" reactiontime="+68" points="563">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Northern Mariana Islands">
              <RESULTS>
                <RESULT eventid="27" place="24" lane="2" heat="4" swimtime="00:01:46.79" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:23.31" />
                    <SPLIT distance="75" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:00:48.51" />
                    <SPLIT distance="125" swimtime="00:01:02.02" />
                    <SPLIT distance="150" swimtime="00:01:16.83" />
                    <SPLIT distance="175" swimtime="00:01:31.19" />
                    <SPLIT distance="200" swimtime="00:01:46.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214457" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="161275" reactiontime="+46" />
                    <RELAYPOSITION number="3" athleteid="201852" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="197310" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Northern Mariana Islands">
              <RESULTS>
                <RESULT eventid="11" place="27" lane="8" heat="2" swimtime="00:01:58.93" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:25.84" />
                    <SPLIT distance="75" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:00:57.47" />
                    <SPLIT distance="125" swimtime="00:01:11.79" />
                    <SPLIT distance="150" swimtime="00:01:29.11" />
                    <SPLIT distance="175" swimtime="00:01:43.29" />
                    <SPLIT distance="200" swimtime="00:01:58.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="214457" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="161275" reactiontime="+41" />
                    <RELAYPOSITION number="3" athleteid="201852" reactiontime="+22" />
                    <RELAYPOSITION number="4" athleteid="197310" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Norway" shortname="NOR" code="NOR" nation="NOR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="130296" lastname="LIE" firstname="Markus" gender="M" birthdate="1995-06-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.00" eventid="3" heat="4" lane="2">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.60" eventid="19" heat="4" lane="7">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:53.03" eventid="23" heat="4" lane="7">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="15" lane="2" heat="4" heatid="40003" swimtime="00:00:50.89" reactiontime="+54" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:24.48" />
                    <SPLIT distance="75" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:00:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="13" lane="8" heat="2" heatid="20203" swimtime="00:00:50.67" reactiontime="+53" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                    <SPLIT distance="50" swimtime="00:00:24.22" />
                    <SPLIT distance="75" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:00:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="22" lane="7" heat="4" heatid="40019" swimtime="00:00:23.65" reactiontime="+54" points="829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:23.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="16" lane="7" heat="4" heatid="40023" swimtime="00:00:52.77" reactiontime="+65" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.90" />
                    <SPLIT distance="50" swimtime="00:00:23.72" />
                    <SPLIT distance="75" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:00:52.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="15" lane="8" heat="1" heatid="10223" swimtime="00:00:52.93" reactiontime="+64" points="807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.54" />
                    <SPLIT distance="50" swimtime="00:00:23.43" />
                    <SPLIT distance="75" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:00:52.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157095" lastname="HAARSAKER" firstname="Christoffer Tofte" gender="M" birthdate="1993-09-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.30" eventid="16" heat="5" lane="3">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.45" eventid="29" heat="3" lane="1">
                  <MEETINFO date="2021-11-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:26.44" eventid="41" heat="8" lane="7">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="33" lane="3" heat="5" heatid="50016" swimtime="00:00:59.13" reactiontime="+70" points="817">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.76" />
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="75" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="22" lane="1" heat="3" heatid="30029" swimtime="00:02:08.80" reactiontime="+76" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="75" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:01.10" />
                    <SPLIT distance="125" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:01:34.60" />
                    <SPLIT distance="175" swimtime="00:01:51.62" />
                    <SPLIT distance="200" swimtime="00:02:08.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="27" lane="7" heat="8" heatid="80041" swimtime="00:00:27.05" reactiontime="+68" points="784">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196342" lastname="LIA" firstname="Nicholas" gender="M" birthdate="2001-02-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.92" eventid="14" heat="8" lane="7">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.56" eventid="5" heat="10" lane="7">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.44" eventid="31" heat="8" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="31" lane="7" heat="8" heatid="80014" swimtime="00:00:47.55" reactiontime="+61" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.75" />
                    <SPLIT distance="50" swimtime="00:00:22.66" />
                    <SPLIT distance="75" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:00:47.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="30" lane="7" heat="10" heatid="100005" swimtime="00:00:23.00" reactiontime="+59" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.35" />
                    <SPLIT distance="50" swimtime="00:00:23.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="27" lane="3" heat="8" heatid="80031" swimtime="00:00:21.43" reactiontime="+59" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:21.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108923" lastname="CHRISTIANSEN" firstname="Henrik" gender="M" birthdate="1996-10-09">
              <ENTRIES>
                <ENTRY entrytime="00:14:30.78" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="00:07:36.57" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="3" lane="2" heat="5" heatid="30110" swimtime="00:14:24.08" reactiontime="+75" points="941">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                    <SPLIT distance="75" swimtime="00:00:40.92" />
                    <SPLIT distance="100" swimtime="00:00:55.32" />
                    <SPLIT distance="125" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:24.48" />
                    <SPLIT distance="175" swimtime="00:01:39.09" />
                    <SPLIT distance="200" swimtime="00:01:53.55" />
                    <SPLIT distance="225" swimtime="00:02:08.10" />
                    <SPLIT distance="250" swimtime="00:02:22.45" />
                    <SPLIT distance="275" swimtime="00:02:36.97" />
                    <SPLIT distance="300" swimtime="00:02:51.31" />
                    <SPLIT distance="325" swimtime="00:03:05.84" />
                    <SPLIT distance="350" swimtime="00:03:20.20" />
                    <SPLIT distance="375" swimtime="00:03:34.63" />
                    <SPLIT distance="400" swimtime="00:03:48.91" />
                    <SPLIT distance="425" swimtime="00:04:03.30" />
                    <SPLIT distance="450" swimtime="00:04:17.49" />
                    <SPLIT distance="475" swimtime="00:04:31.89" />
                    <SPLIT distance="500" swimtime="00:04:46.09" />
                    <SPLIT distance="525" swimtime="00:05:00.38" />
                    <SPLIT distance="550" swimtime="00:05:14.68" />
                    <SPLIT distance="575" swimtime="00:05:28.98" />
                    <SPLIT distance="600" swimtime="00:05:43.29" />
                    <SPLIT distance="625" swimtime="00:05:57.48" />
                    <SPLIT distance="650" swimtime="00:06:11.78" />
                    <SPLIT distance="675" swimtime="00:06:26.09" />
                    <SPLIT distance="700" swimtime="00:06:40.34" />
                    <SPLIT distance="725" swimtime="00:06:54.56" />
                    <SPLIT distance="750" swimtime="00:07:08.72" />
                    <SPLIT distance="775" swimtime="00:07:23.00" />
                    <SPLIT distance="800" swimtime="00:07:37.35" />
                    <SPLIT distance="825" swimtime="00:07:51.61" />
                    <SPLIT distance="850" swimtime="00:08:05.79" />
                    <SPLIT distance="875" swimtime="00:08:20.05" />
                    <SPLIT distance="900" swimtime="00:08:34.14" />
                    <SPLIT distance="925" swimtime="00:08:48.38" />
                    <SPLIT distance="950" swimtime="00:09:02.56" />
                    <SPLIT distance="975" swimtime="00:09:16.67" />
                    <SPLIT distance="1000" swimtime="00:09:30.93" />
                    <SPLIT distance="1025" swimtime="00:09:45.29" />
                    <SPLIT distance="1050" swimtime="00:09:59.62" />
                    <SPLIT distance="1075" swimtime="00:10:14.04" />
                    <SPLIT distance="1100" swimtime="00:10:28.24" />
                    <SPLIT distance="1125" swimtime="00:10:42.70" />
                    <SPLIT distance="1150" swimtime="00:10:57.04" />
                    <SPLIT distance="1175" swimtime="00:11:11.74" />
                    <SPLIT distance="1200" swimtime="00:11:26.33" />
                    <SPLIT distance="1225" swimtime="00:11:40.87" />
                    <SPLIT distance="1250" swimtime="00:11:55.41" />
                    <SPLIT distance="1275" swimtime="00:12:10.05" />
                    <SPLIT distance="1300" swimtime="00:12:24.67" />
                    <SPLIT distance="1325" swimtime="00:12:39.36" />
                    <SPLIT distance="1350" swimtime="00:12:54.17" />
                    <SPLIT distance="1375" swimtime="00:13:09.10" />
                    <SPLIT distance="1400" swimtime="00:13:24.29" />
                    <SPLIT distance="1425" swimtime="00:13:39.67" />
                    <SPLIT distance="1450" swimtime="00:13:54.97" />
                    <SPLIT distance="1475" swimtime="00:14:10.02" />
                    <SPLIT distance="1500" swimtime="00:14:24.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="2" lane="2" heat="5" heatid="30142" swimtime="00:07:31.48" reactiontime="+74" points="947">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="75" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:00:55.35" />
                    <SPLIT distance="125" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:24.03" />
                    <SPLIT distance="175" swimtime="00:01:38.36" />
                    <SPLIT distance="200" swimtime="00:01:52.73" />
                    <SPLIT distance="225" swimtime="00:02:07.07" />
                    <SPLIT distance="250" swimtime="00:02:21.24" />
                    <SPLIT distance="275" swimtime="00:02:35.36" />
                    <SPLIT distance="300" swimtime="00:02:49.60" />
                    <SPLIT distance="325" swimtime="00:03:03.87" />
                    <SPLIT distance="350" swimtime="00:03:18.06" />
                    <SPLIT distance="375" swimtime="00:03:32.34" />
                    <SPLIT distance="400" swimtime="00:03:46.52" />
                    <SPLIT distance="425" swimtime="00:04:00.74" />
                    <SPLIT distance="450" swimtime="00:04:14.94" />
                    <SPLIT distance="475" swimtime="00:04:29.05" />
                    <SPLIT distance="500" swimtime="00:04:43.18" />
                    <SPLIT distance="525" swimtime="00:04:57.23" />
                    <SPLIT distance="550" swimtime="00:05:11.47" />
                    <SPLIT distance="575" swimtime="00:05:25.55" />
                    <SPLIT distance="600" swimtime="00:05:39.57" />
                    <SPLIT distance="625" swimtime="00:05:53.61" />
                    <SPLIT distance="650" swimtime="00:06:07.66" />
                    <SPLIT distance="675" swimtime="00:06:21.67" />
                    <SPLIT distance="700" swimtime="00:06:35.92" />
                    <SPLIT distance="725" swimtime="00:06:49.93" />
                    <SPLIT distance="750" swimtime="00:07:04.09" />
                    <SPLIT distance="775" swimtime="00:07:17.83" />
                    <SPLIT distance="800" swimtime="00:07:31.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197436" lastname="JOENTVEDT" firstname="Jon" gender="M" birthdate="2003-07-28">
              <ENTRIES>
                <ENTRY entrytime="00:14:45.19" eventid="10" heat="2" lane="6">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:03:43.24" eventid="24" heat="3" lane="5">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="35" />
                <ENTRY entrytime="00:07:52.21" eventid="42" heat="1" lane="4">
                  <MEETINFO date="2022-04-01" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="-1" lane="6" heat="2" heatid="20010" swimtime="NT" status="DNS" />
                <RESULT eventid="24" place="-1" lane="5" heat="3" heatid="30024" swimtime="NT" status="DNS" />
                <RESULT eventid="142" place="18" lane="4" heat="1" heatid="10042" swimtime="00:07:55.93" reactiontime="+73" points="808">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                    <SPLIT distance="75" swimtime="00:00:41.03" />
                    <SPLIT distance="100" swimtime="00:00:55.47" />
                    <SPLIT distance="125" swimtime="00:01:10.10" />
                    <SPLIT distance="150" swimtime="00:01:24.67" />
                    <SPLIT distance="175" swimtime="00:01:39.37" />
                    <SPLIT distance="200" swimtime="00:01:54.06" />
                    <SPLIT distance="225" swimtime="00:02:09.25" />
                    <SPLIT distance="250" swimtime="00:02:24.11" />
                    <SPLIT distance="275" swimtime="00:02:39.07" />
                    <SPLIT distance="300" swimtime="00:02:54.20" />
                    <SPLIT distance="325" swimtime="00:03:09.26" />
                    <SPLIT distance="350" swimtime="00:03:24.63" />
                    <SPLIT distance="375" swimtime="00:03:40.03" />
                    <SPLIT distance="400" swimtime="00:03:55.31" />
                    <SPLIT distance="425" swimtime="00:04:10.55" />
                    <SPLIT distance="450" swimtime="00:04:25.95" />
                    <SPLIT distance="475" swimtime="00:04:41.33" />
                    <SPLIT distance="500" swimtime="00:04:56.66" />
                    <SPLIT distance="525" swimtime="00:05:11.99" />
                    <SPLIT distance="550" swimtime="00:05:27.24" />
                    <SPLIT distance="575" swimtime="00:05:42.08" />
                    <SPLIT distance="600" swimtime="00:05:57.34" />
                    <SPLIT distance="625" swimtime="00:06:12.47" />
                    <SPLIT distance="650" swimtime="00:06:27.67" />
                    <SPLIT distance="675" swimtime="00:06:42.86" />
                    <SPLIT distance="700" swimtime="00:06:57.94" />
                    <SPLIT distance="725" swimtime="00:07:13.05" />
                    <SPLIT distance="750" swimtime="00:07:28.29" />
                    <SPLIT distance="775" swimtime="00:07:42.42" />
                    <SPLIT distance="800" swimtime="00:07:55.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157016" lastname="LØYNING" firstname="Ingeborg" gender="F" birthdate="2000-09-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.15" eventid="2" heat="5" lane="2">
                  <MEETINFO date="2021-09-25" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.67" eventid="45" heat="3" lane="3">
                  <MEETINFO date="2021-09-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.47" eventid="18" heat="5" lane="2">
                  <MEETINFO date="2021-09-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="23" lane="2" heat="5" heatid="50002" swimtime="00:00:58.49" reactiontime="+59" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                    <SPLIT distance="75" swimtime="00:00:43.21" />
                    <SPLIT distance="100" swimtime="00:00:58.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="22" lane="3" heat="3" heatid="30045" swimtime="00:02:07.67" reactiontime="+55" points="808">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.06" />
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="75" swimtime="00:00:44.75" />
                    <SPLIT distance="100" swimtime="00:01:00.40" />
                    <SPLIT distance="125" swimtime="00:01:16.52" />
                    <SPLIT distance="150" swimtime="00:01:33.06" />
                    <SPLIT distance="175" swimtime="00:01:50.11" />
                    <SPLIT distance="200" swimtime="00:02:07.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="25" lane="2" heat="5" heatid="50018" swimtime="00:00:27.20" reactiontime="+55" points="801">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212842" lastname="SLYNGSTADLI" firstname="Silje" gender="F" birthdate="2004-04-01">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.88" eventid="15" heat="4" lane="1">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.34" eventid="40" heat="5" lane="1">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="-1" lane="1" heat="4" heatid="40015" swimtime="NT" status="DNS" />
                <RESULT eventid="40" place="18" lane="1" heat="5" heatid="50040" swimtime="00:00:30.36" reactiontime="+66" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Norway">
              <RESULTS>
                <RESULT eventid="48" place="12" lane="5" heat="2" swimtime="00:03:28.97" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:24.71" />
                    <SPLIT distance="75" swimtime="00:00:37.75" />
                    <SPLIT distance="100" swimtime="00:00:50.76" />
                    <SPLIT distance="125" swimtime="00:01:02.76" />
                    <SPLIT distance="150" swimtime="00:01:17.84" />
                    <SPLIT distance="175" swimtime="00:01:33.14" />
                    <SPLIT distance="200" swimtime="00:01:48.87" />
                    <SPLIT distance="225" swimtime="00:01:59.81" />
                    <SPLIT distance="250" swimtime="00:02:13.22" />
                    <SPLIT distance="275" swimtime="00:02:27.42" />
                    <SPLIT distance="300" swimtime="00:02:42.45" />
                    <SPLIT distance="325" swimtime="00:02:52.66" />
                    <SPLIT distance="350" swimtime="00:03:04.57" />
                    <SPLIT distance="375" swimtime="00:03:16.90" />
                    <SPLIT distance="400" swimtime="00:03:28.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130296" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="157095" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="197436" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="196342" reactiontime="+9" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Norway">
              <RESULTS>
                <RESULT eventid="35" place="10" lane="2" heat="3" swimtime="00:01:34.43" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:23.62" />
                    <SPLIT distance="75" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:00:49.97" />
                    <SPLIT distance="125" swimtime="00:01:00.64" />
                    <SPLIT distance="150" swimtime="00:01:13.74" />
                    <SPLIT distance="175" swimtime="00:01:23.35" />
                    <SPLIT distance="200" swimtime="00:01:34.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="130296" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="157095" reactiontime="+10" />
                    <RELAYPOSITION number="3" athleteid="197436" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="196342" reactiontime="+6" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="New Zealand" shortname="NZL" code="NZL" nation="NZL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="161935" lastname="DELL" firstname="Zac" gender="M" birthdate="2001-01-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.61" eventid="3" heat="6" lane="1">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="24" lane="1" heat="6" heatid="60003" swimtime="00:00:51.98" reactiontime="+56" points="803">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:24.64" />
                    <SPLIT distance="75" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:00:51.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212856" lastname="GILBERT" firstname="Josh" gender="M" birthdate="2001-06-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.33" eventid="16" heat="4" lane="7">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.27" eventid="29" heat="4" lane="8">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:27.05" eventid="41" heat="6" lane="7">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="21" lane="7" heat="4" heatid="40016" swimtime="00:00:58.06" reactiontime="+62" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:26.99" />
                    <SPLIT distance="75" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:00:58.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="20" lane="8" heat="4" heatid="40029" swimtime="00:02:08.27" reactiontime="+63" points="822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                    <SPLIT distance="75" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:01.73" />
                    <SPLIT distance="125" swimtime="00:01:18.21" />
                    <SPLIT distance="150" swimtime="00:01:34.91" />
                    <SPLIT distance="175" swimtime="00:01:51.34" />
                    <SPLIT distance="200" swimtime="00:02:08.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="25" lane="7" heat="6" heatid="60041" swimtime="00:00:26.95" reactiontime="+61" points="793">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202034" lastname="GRAY" firstname="Cameron" gender="M" birthdate="2003-08-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.58" eventid="39" heat="5" lane="8">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.74" eventid="19" heat="5" lane="8">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.05" eventid="5" heat="7" lane="6">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.76" eventid="31" heat="8" lane="7">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="26" lane="8" heat="5" heatid="50039" swimtime="00:00:51.69" reactiontime="+67" points="789">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.97" />
                    <SPLIT distance="50" swimtime="00:00:24.03" />
                    <SPLIT distance="75" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="18" lane="8" heat="5" heatid="50019" swimtime="00:00:23.49" reactiontime="+61" points="846">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:23.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="26" lane="6" heat="7" heatid="70005" swimtime="00:00:22.90" reactiontime="+68" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.51" />
                    <SPLIT distance="50" swimtime="00:00:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="30" lane="7" heat="8" heatid="80031" swimtime="00:00:21.50" reactiontime="+67" points="824">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.35" />
                    <SPLIT distance="50" swimtime="00:00:21.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202035" lastname="SWIFT" firstname="Carter" gender="M" birthdate="1998-12-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.17" eventid="14" heat="9" lane="8">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.49" eventid="44" heat="4" lane="8">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="27" lane="8" heat="9" heatid="90014" swimtime="00:00:47.36" reactiontime="+62" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.54" />
                    <SPLIT distance="75" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:00:47.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="22" lane="8" heat="4" heatid="40044" swimtime="00:01:44.88" reactiontime="+60" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.30" />
                    <SPLIT distance="50" swimtime="00:00:24.19" />
                    <SPLIT distance="75" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:00:50.45" />
                    <SPLIT distance="125" swimtime="00:01:03.94" />
                    <SPLIT distance="150" swimtime="00:01:17.51" />
                    <SPLIT distance="175" swimtime="00:01:31.27" />
                    <SPLIT distance="200" swimtime="00:01:44.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212853" lastname="FOLLOWS" firstname="Kane" gender="M" birthdate="1997-05-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.05" eventid="46" heat="3" lane="1">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="14" lane="1" heat="3" heatid="30046" swimtime="00:01:53.11" reactiontime="+62" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.70" />
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                    <SPLIT distance="75" swimtime="00:00:40.68" />
                    <SPLIT distance="100" swimtime="00:00:54.81" />
                    <SPLIT distance="125" swimtime="00:01:08.96" />
                    <SPLIT distance="150" swimtime="00:01:23.42" />
                    <SPLIT distance="175" swimtime="00:01:38.33" />
                    <SPLIT distance="200" swimtime="00:01:53.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="162436" lastname="GROBBELAAR" firstname="Luan" gender="M" birthdate="2002-03-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:57.77" eventid="7" heat="2" lane="4">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="00:04:10.47" eventid="37" heat="2" lane="8">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="23" lane="4" heat="2" heatid="20007" swimtime="00:01:57.38" reactiontime="+67" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:00:55.82" />
                    <SPLIT distance="125" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:29.26" />
                    <SPLIT distance="175" swimtime="00:01:43.88" />
                    <SPLIT distance="200" swimtime="00:01:57.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="13" lane="8" heat="2" heatid="20037" swimtime="00:04:09.98" reactiontime="+67" points="828">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="75" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:00:57.42" />
                    <SPLIT distance="125" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:29.41" />
                    <SPLIT distance="175" swimtime="00:01:44.93" />
                    <SPLIT distance="200" swimtime="00:02:00.45" />
                    <SPLIT distance="225" swimtime="00:02:17.97" />
                    <SPLIT distance="250" swimtime="00:02:35.48" />
                    <SPLIT distance="275" swimtime="00:02:53.25" />
                    <SPLIT distance="300" swimtime="00:03:11.08" />
                    <SPLIT distance="325" swimtime="00:03:26.53" />
                    <SPLIT distance="350" swimtime="00:03:41.09" />
                    <SPLIT distance="375" swimtime="00:03:55.78" />
                    <SPLIT distance="400" swimtime="00:04:09.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164930" lastname="CLARK" firstname="Louis" gender="M" birthdate="2001-08-21">
              <ENTRIES>
                <ENTRY entrytime="00:03:45.94" eventid="24" heat="3" lane="2">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="00:07:49.54" eventid="42" heat="2" lane="6">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="24" place="20" lane="2" heat="3" heatid="30024" swimtime="00:03:46.19" reactiontime="+76" points="826">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:25.52" />
                    <SPLIT distance="75" swimtime="00:00:39.44" />
                    <SPLIT distance="100" swimtime="00:00:53.61" />
                    <SPLIT distance="125" swimtime="00:01:07.62" />
                    <SPLIT distance="150" swimtime="00:01:21.93" />
                    <SPLIT distance="175" swimtime="00:01:36.34" />
                    <SPLIT distance="200" swimtime="00:01:50.71" />
                    <SPLIT distance="225" swimtime="00:02:05.10" />
                    <SPLIT distance="250" swimtime="00:02:19.52" />
                    <SPLIT distance="275" swimtime="00:02:34.05" />
                    <SPLIT distance="300" swimtime="00:02:48.60" />
                    <SPLIT distance="325" swimtime="00:03:02.95" />
                    <SPLIT distance="350" swimtime="00:03:17.67" />
                    <SPLIT distance="375" swimtime="00:03:32.10" />
                    <SPLIT distance="400" swimtime="00:03:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="16" lane="6" heat="2" heatid="20042" swimtime="00:07:53.36" reactiontime="+69" points="821">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="75" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:00:55.39" />
                    <SPLIT distance="125" swimtime="00:01:09.99" />
                    <SPLIT distance="150" swimtime="00:01:24.73" />
                    <SPLIT distance="175" swimtime="00:01:39.42" />
                    <SPLIT distance="200" swimtime="00:01:54.10" />
                    <SPLIT distance="225" swimtime="00:02:08.51" />
                    <SPLIT distance="250" swimtime="00:02:23.17" />
                    <SPLIT distance="275" swimtime="00:02:37.72" />
                    <SPLIT distance="300" swimtime="00:02:52.39" />
                    <SPLIT distance="325" swimtime="00:03:07.02" />
                    <SPLIT distance="350" swimtime="00:03:21.76" />
                    <SPLIT distance="375" swimtime="00:03:36.53" />
                    <SPLIT distance="400" swimtime="00:03:51.50" />
                    <SPLIT distance="425" swimtime="00:04:06.53" />
                    <SPLIT distance="450" swimtime="00:04:21.49" />
                    <SPLIT distance="475" swimtime="00:04:36.30" />
                    <SPLIT distance="500" swimtime="00:04:51.53" />
                    <SPLIT distance="525" swimtime="00:05:06.55" />
                    <SPLIT distance="550" swimtime="00:05:21.69" />
                    <SPLIT distance="575" swimtime="00:05:36.64" />
                    <SPLIT distance="600" swimtime="00:05:51.90" />
                    <SPLIT distance="625" swimtime="00:06:07.09" />
                    <SPLIT distance="650" swimtime="00:06:22.21" />
                    <SPLIT distance="675" swimtime="00:06:37.35" />
                    <SPLIT distance="700" swimtime="00:06:52.65" />
                    <SPLIT distance="725" swimtime="00:07:07.96" />
                    <SPLIT distance="750" swimtime="00:07:23.45" />
                    <SPLIT distance="775" swimtime="00:07:38.81" />
                    <SPLIT distance="800" swimtime="00:07:53.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156844" lastname="OUWEHAND" firstname="Vanessa Hazel" gender="F" birthdate="1999-12-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.31" eventid="2" heat="3" lane="5">
                  <MEETINFO date="2021-08-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="25" lane="5" heat="3" heatid="30002" swimtime="00:00:58.56" reactiontime="+57" points="823">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                    <SPLIT distance="75" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:00:58.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143885" lastname="GASSON" firstname="Helena" gender="F" birthdate="1994-12-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.04" eventid="38" heat="4" lane="2">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.39" eventid="6" heat="5" lane="2">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.50" eventid="4" heat="5" lane="2">
                  <MEETINFO date="2021-08-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.78" eventid="22" heat="4" lane="3">
                  <MEETINFO date="2021-08-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="15" lane="2" heat="4" heatid="40038" swimtime="00:00:57.51" reactiontime="+60" points="855">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                    <SPLIT distance="75" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="14" lane="8" heat="2" heatid="20238" swimtime="00:00:57.23" reactiontime="+63" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="75" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:00:57.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="19" lane="2" heat="5" heatid="50006" swimtime="00:02:10.33" reactiontime="+63" points="817">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.28" />
                    <SPLIT distance="50" swimtime="00:00:27.56" />
                    <SPLIT distance="75" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:00.41" />
                    <SPLIT distance="125" swimtime="00:01:19.08" />
                    <SPLIT distance="150" swimtime="00:01:38.55" />
                    <SPLIT distance="175" swimtime="00:01:55.31" />
                    <SPLIT distance="200" swimtime="00:02:10.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="15" lane="2" heat="5" heatid="50004" swimtime="00:00:25.63" reactiontime="+63" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:25.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="11" lane="8" heat="2" heatid="20204" swimtime="00:00:25.38" reactiontime="+63" points="886">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="5" lane="8" heat="1" heatid="10122" swimtime="00:00:58.40" reactiontime="+61" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                    <SPLIT distance="75" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:00:58.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="3" lane="3" heat="4" heatid="40022" swimtime="00:00:58.92" reactiontime="+61" points="882">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:26.51" />
                    <SPLIT distance="75" swimtime="00:00:43.67" />
                    <SPLIT distance="100" swimtime="00:00:58.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="8" lane="5" heat="2" heatid="20222" swimtime="00:00:59.15" reactiontime="+63" points="871">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:26.25" />
                    <SPLIT distance="75" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:00:59.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156788" lastname="GODWIN" firstname="Emma" gender="F" birthdate="1997-04-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:02:07.11" eventid="45" heat="4" lane="1">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:27.35" eventid="18" heat="5" lane="1">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="23" lane="1" heat="4" heatid="40045" swimtime="00:02:07.91" reactiontime="+57" points="804">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="75" swimtime="00:00:45.93" />
                    <SPLIT distance="100" swimtime="00:01:02.19" />
                    <SPLIT distance="125" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:01:34.70" />
                    <SPLIT distance="175" swimtime="00:01:51.29" />
                    <SPLIT distance="200" swimtime="00:02:07.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="28" lane="1" heat="5" heatid="50018" swimtime="00:00:27.37" reactiontime="+58" points="787">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212855" lastname="PATERSON" firstname="Esme" gender="F" birthdate="2001-09-24">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.99" eventid="20" heat="1" lane="4">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="-1" lane="4" heat="1" heatid="10020" swimtime="00:02:11.75" status="DSQ" reactiontime="+72" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156786" lastname="DEANS" firstname="Caitlin" gender="F" birthdate="1999-12-05">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.10" eventid="43" heat="3" lane="8">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:16:05.52" eventid="33" heat="0" lane="-1">
                  <MEETINFO date="2022-08-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="19" lane="8" heat="3" heatid="30043" swimtime="00:01:57.93" reactiontime="+75" points="818">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.47" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="75" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:00:57.57" />
                    <SPLIT distance="125" swimtime="00:01:12.67" />
                    <SPLIT distance="150" swimtime="00:01:27.67" />
                    <SPLIT distance="175" swimtime="00:01:43.06" />
                    <SPLIT distance="200" swimtime="00:01:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="5" lane="1" heat="5" heatid="30133" swimtime="00:15:51.98" reactiontime="+77" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                    <SPLIT distance="75" swimtime="00:00:44.22" />
                    <SPLIT distance="100" swimtime="00:00:59.81" />
                    <SPLIT distance="125" swimtime="00:01:15.66" />
                    <SPLIT distance="150" swimtime="00:01:31.69" />
                    <SPLIT distance="175" swimtime="00:01:47.72" />
                    <SPLIT distance="200" swimtime="00:02:03.72" />
                    <SPLIT distance="225" swimtime="00:02:19.67" />
                    <SPLIT distance="250" swimtime="00:02:35.63" />
                    <SPLIT distance="275" swimtime="00:02:51.60" />
                    <SPLIT distance="300" swimtime="00:03:07.45" />
                    <SPLIT distance="325" swimtime="00:03:23.33" />
                    <SPLIT distance="350" swimtime="00:03:39.19" />
                    <SPLIT distance="375" swimtime="00:03:54.96" />
                    <SPLIT distance="400" swimtime="00:04:10.82" />
                    <SPLIT distance="425" swimtime="00:04:26.59" />
                    <SPLIT distance="450" swimtime="00:04:42.53" />
                    <SPLIT distance="475" swimtime="00:04:58.40" />
                    <SPLIT distance="500" swimtime="00:05:14.46" />
                    <SPLIT distance="525" swimtime="00:05:30.32" />
                    <SPLIT distance="550" swimtime="00:05:46.35" />
                    <SPLIT distance="575" swimtime="00:06:02.17" />
                    <SPLIT distance="600" swimtime="00:06:18.10" />
                    <SPLIT distance="625" swimtime="00:06:34.19" />
                    <SPLIT distance="650" swimtime="00:06:50.15" />
                    <SPLIT distance="675" swimtime="00:07:06.14" />
                    <SPLIT distance="700" swimtime="00:07:22.15" />
                    <SPLIT distance="725" swimtime="00:07:38.10" />
                    <SPLIT distance="750" swimtime="00:07:54.06" />
                    <SPLIT distance="775" swimtime="00:08:10.08" />
                    <SPLIT distance="800" swimtime="00:08:26.14" />
                    <SPLIT distance="825" swimtime="00:08:42.06" />
                    <SPLIT distance="850" swimtime="00:08:58.06" />
                    <SPLIT distance="875" swimtime="00:09:13.92" />
                    <SPLIT distance="900" swimtime="00:09:29.80" />
                    <SPLIT distance="925" swimtime="00:09:45.68" />
                    <SPLIT distance="950" swimtime="00:10:01.75" />
                    <SPLIT distance="975" swimtime="00:10:17.70" />
                    <SPLIT distance="1000" swimtime="00:10:33.61" />
                    <SPLIT distance="1025" swimtime="00:10:49.59" />
                    <SPLIT distance="1050" swimtime="00:11:05.67" />
                    <SPLIT distance="1075" swimtime="00:11:21.70" />
                    <SPLIT distance="1100" swimtime="00:11:37.73" />
                    <SPLIT distance="1125" swimtime="00:11:53.63" />
                    <SPLIT distance="1150" swimtime="00:12:09.69" />
                    <SPLIT distance="1175" swimtime="00:12:25.57" />
                    <SPLIT distance="1200" swimtime="00:12:41.49" />
                    <SPLIT distance="1225" swimtime="00:12:57.57" />
                    <SPLIT distance="1250" swimtime="00:13:13.68" />
                    <SPLIT distance="1275" swimtime="00:13:29.74" />
                    <SPLIT distance="1300" swimtime="00:13:45.94" />
                    <SPLIT distance="1325" swimtime="00:14:02.12" />
                    <SPLIT distance="1350" swimtime="00:14:18.23" />
                    <SPLIT distance="1375" swimtime="00:14:34.43" />
                    <SPLIT distance="1400" swimtime="00:14:50.46" />
                    <SPLIT distance="1425" swimtime="00:15:06.28" />
                    <SPLIT distance="1450" swimtime="00:15:21.89" />
                    <SPLIT distance="1475" swimtime="00:15:37.12" />
                    <SPLIT distance="1500" swimtime="00:15:51.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161792" lastname="FAIRWEATHER" firstname="Erika" gender="F" birthdate="2003-12-31">
              <ENTRIES>
                <ENTRY entrytime="00:04:02.28" eventid="1" heat="4" lane="2">
                  <MEETINFO date="2021-07-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:08:18.63" eventid="12" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="101" place="2" lane="4" heat="1" heatid="10101" swimtime="00:03:56.00" reactiontime="+70" points="973">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.75" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:41.72" />
                    <SPLIT distance="100" swimtime="00:00:56.59" />
                    <SPLIT distance="125" swimtime="00:01:11.53" />
                    <SPLIT distance="150" swimtime="00:01:26.59" />
                    <SPLIT distance="175" swimtime="00:01:41.62" />
                    <SPLIT distance="200" swimtime="00:01:56.69" />
                    <SPLIT distance="225" swimtime="00:02:11.57" />
                    <SPLIT distance="250" swimtime="00:02:26.61" />
                    <SPLIT distance="275" swimtime="00:02:41.64" />
                    <SPLIT distance="300" swimtime="00:02:56.67" />
                    <SPLIT distance="325" swimtime="00:03:11.77" />
                    <SPLIT distance="350" swimtime="00:03:26.75" />
                    <SPLIT distance="375" swimtime="00:03:41.77" />
                    <SPLIT distance="400" swimtime="00:03:56.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="1" lane="2" heat="4" heatid="40001" swimtime="00:03:58.27" reactiontime="+72" points="946">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="75" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:00:56.78" />
                    <SPLIT distance="125" swimtime="00:01:11.77" />
                    <SPLIT distance="150" swimtime="00:01:26.90" />
                    <SPLIT distance="175" swimtime="00:01:41.96" />
                    <SPLIT distance="200" swimtime="00:01:57.14" />
                    <SPLIT distance="225" swimtime="00:02:12.18" />
                    <SPLIT distance="250" swimtime="00:02:27.42" />
                    <SPLIT distance="275" swimtime="00:02:42.63" />
                    <SPLIT distance="300" swimtime="00:02:57.99" />
                    <SPLIT distance="325" swimtime="00:03:13.27" />
                    <SPLIT distance="350" swimtime="00:03:28.56" />
                    <SPLIT distance="375" swimtime="00:03:43.70" />
                    <SPLIT distance="400" swimtime="00:03:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="2" lane="7" heat="5" heatid="30112" swimtime="00:08:10.41" reactiontime="+72" points="933">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="75" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:00:58.36" />
                    <SPLIT distance="125" swimtime="00:01:13.66" />
                    <SPLIT distance="150" swimtime="00:01:29.06" />
                    <SPLIT distance="175" swimtime="00:01:44.29" />
                    <SPLIT distance="200" swimtime="00:01:59.69" />
                    <SPLIT distance="225" swimtime="00:02:15.00" />
                    <SPLIT distance="250" swimtime="00:02:30.49" />
                    <SPLIT distance="275" swimtime="00:02:45.99" />
                    <SPLIT distance="300" swimtime="00:03:01.49" />
                    <SPLIT distance="325" swimtime="00:03:16.86" />
                    <SPLIT distance="350" swimtime="00:03:32.41" />
                    <SPLIT distance="375" swimtime="00:03:47.76" />
                    <SPLIT distance="400" swimtime="00:04:03.22" />
                    <SPLIT distance="425" swimtime="00:04:18.69" />
                    <SPLIT distance="450" swimtime="00:04:34.21" />
                    <SPLIT distance="475" swimtime="00:04:49.68" />
                    <SPLIT distance="500" swimtime="00:05:05.37" />
                    <SPLIT distance="525" swimtime="00:05:21.02" />
                    <SPLIT distance="550" swimtime="00:05:36.80" />
                    <SPLIT distance="575" swimtime="00:05:52.30" />
                    <SPLIT distance="600" swimtime="00:06:07.95" />
                    <SPLIT distance="625" swimtime="00:06:23.59" />
                    <SPLIT distance="650" swimtime="00:06:39.42" />
                    <SPLIT distance="675" swimtime="00:06:54.81" />
                    <SPLIT distance="700" swimtime="00:07:10.39" />
                    <SPLIT distance="725" swimtime="00:07:25.86" />
                    <SPLIT distance="750" swimtime="00:07:41.60" />
                    <SPLIT distance="775" swimtime="00:07:56.24" />
                    <SPLIT distance="800" swimtime="00:08:10.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201331" lastname="RASMUSSEN" firstname="Mya" gender="F" birthdate="2000-06-21">
              <ENTRIES>
                <ENTRY entrytime="00:04:41.81" eventid="36" heat="2" lane="2">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="36" place="12" lane="2" heat="2" heatid="20036" swimtime="00:04:36.08" reactiontime="+58" points="825">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.85" />
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="75" swimtime="00:00:46.68" />
                    <SPLIT distance="100" swimtime="00:01:03.65" />
                    <SPLIT distance="125" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:01:39.00" />
                    <SPLIT distance="175" swimtime="00:01:56.62" />
                    <SPLIT distance="200" swimtime="00:02:14.35" />
                    <SPLIT distance="225" swimtime="00:02:33.48" />
                    <SPLIT distance="250" swimtime="00:02:52.90" />
                    <SPLIT distance="275" swimtime="00:03:12.21" />
                    <SPLIT distance="300" swimtime="00:03:31.89" />
                    <SPLIT distance="325" swimtime="00:03:48.50" />
                    <SPLIT distance="350" swimtime="00:04:04.45" />
                    <SPLIT distance="375" swimtime="00:04:20.47" />
                    <SPLIT distance="400" swimtime="00:04:36.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156796" lastname="MOYNIHAN" firstname="Rebecca" gender="F" birthdate="1998-05-26">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:24.93" eventid="30" heat="6" lane="1">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="30" place="15" lane="1" heat="6" heatid="60030" swimtime="00:00:24.59" reactiontime="+69" points="810">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:24.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="16" lane="8" heat="2" heatid="20230" swimtime="00:00:24.67" reactiontime="+70" points="802">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:24.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214488" lastname="WILLIAMS" firstname="George" gender="M" birthdate="1999-04-17" />
            <ATHLETE athleteid="212851" lastname="LITTLEJOHN" firstname="Ben Jago" gender="M" birthdate="2002-04-03" />
            <ATHLETE athleteid="212854" lastname="OSBORNE" firstname="Summer" gender="F" birthdate="2005-05-23" />
            <ATHLETE athleteid="202036" lastname="HEATH" firstname="Ruby" gender="F" birthdate="1999-12-06" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="New Zealand">
              <RESULTS>
                <RESULT eventid="9" place="9" lane="7" heat="1" swimtime="00:03:10.97" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.60" />
                    <SPLIT distance="50" swimtime="00:00:22.94" />
                    <SPLIT distance="75" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:00:47.93" />
                    <SPLIT distance="125" swimtime="00:00:58.10" />
                    <SPLIT distance="150" swimtime="00:01:10.04" />
                    <SPLIT distance="175" swimtime="00:01:22.37" />
                    <SPLIT distance="200" swimtime="00:01:34.85" />
                    <SPLIT distance="225" swimtime="00:01:45.01" />
                    <SPLIT distance="250" swimtime="00:01:57.02" />
                    <SPLIT distance="275" swimtime="00:02:09.57" />
                    <SPLIT distance="300" swimtime="00:02:22.44" />
                    <SPLIT distance="325" swimtime="00:02:33.35" />
                    <SPLIT distance="350" swimtime="00:02:45.54" />
                    <SPLIT distance="375" swimtime="00:02:58.28" />
                    <SPLIT distance="400" swimtime="00:03:10.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202034" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="202035" reactiontime="+14" />
                    <RELAYPOSITION number="3" athleteid="161935" reactiontime="+21" />
                    <RELAYPOSITION number="4" athleteid="214488" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="New Zealand">
              <RESULTS>
                <RESULT eventid="48" place="10" lane="3" heat="1" swimtime="00:03:26.68" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                    <SPLIT distance="75" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:00:52.19" />
                    <SPLIT distance="125" swimtime="00:01:04.02" />
                    <SPLIT distance="150" swimtime="00:01:18.87" />
                    <SPLIT distance="175" swimtime="00:01:34.44" />
                    <SPLIT distance="200" swimtime="00:01:50.02" />
                    <SPLIT distance="225" swimtime="00:02:00.18" />
                    <SPLIT distance="250" swimtime="00:02:12.99" />
                    <SPLIT distance="275" swimtime="00:02:26.54" />
                    <SPLIT distance="300" swimtime="00:02:40.42" />
                    <SPLIT distance="325" swimtime="00:02:50.57" />
                    <SPLIT distance="350" swimtime="00:03:02.16" />
                    <SPLIT distance="375" swimtime="00:03:14.46" />
                    <SPLIT distance="400" swimtime="00:03:26.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="161935" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="212856" reactiontime="+11" />
                    <RELAYPOSITION number="3" athleteid="202034" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="202035" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="New Zealand">
              <RESULTS>
                <RESULT eventid="32" place="10" lane="7" heat="1" swimtime="00:07:03.11" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                    <SPLIT distance="50" swimtime="00:00:24.31" />
                    <SPLIT distance="75" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:00:50.74" />
                    <SPLIT distance="125" swimtime="00:01:03.90" />
                    <SPLIT distance="150" swimtime="00:01:17.52" />
                    <SPLIT distance="175" swimtime="00:01:31.27" />
                    <SPLIT distance="200" swimtime="00:01:44.60" />
                    <SPLIT distance="225" swimtime="00:01:55.53" />
                    <SPLIT distance="250" swimtime="00:02:08.51" />
                    <SPLIT distance="275" swimtime="00:02:21.91" />
                    <SPLIT distance="300" swimtime="00:02:35.51" />
                    <SPLIT distance="325" swimtime="00:02:49.21" />
                    <SPLIT distance="350" swimtime="00:03:03.01" />
                    <SPLIT distance="375" swimtime="00:03:16.78" />
                    <SPLIT distance="400" swimtime="00:03:30.28" />
                    <SPLIT distance="425" swimtime="00:03:41.20" />
                    <SPLIT distance="450" swimtime="00:03:54.39" />
                    <SPLIT distance="475" swimtime="00:04:07.79" />
                    <SPLIT distance="500" swimtime="00:04:21.27" />
                    <SPLIT distance="525" swimtime="00:04:34.92" />
                    <SPLIT distance="550" swimtime="00:04:48.91" />
                    <SPLIT distance="575" swimtime="00:05:02.99" />
                    <SPLIT distance="600" swimtime="00:05:16.35" />
                    <SPLIT distance="625" swimtime="00:05:27.35" />
                    <SPLIT distance="650" swimtime="00:05:40.37" />
                    <SPLIT distance="675" swimtime="00:05:53.49" />
                    <SPLIT distance="700" swimtime="00:06:06.95" />
                    <SPLIT distance="725" swimtime="00:06:20.60" />
                    <SPLIT distance="750" swimtime="00:06:34.65" />
                    <SPLIT distance="775" swimtime="00:06:49.05" />
                    <SPLIT distance="800" swimtime="00:07:03.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="212851" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="202035" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="202034" reactiontime="+10" />
                    <RELAYPOSITION number="4" athleteid="164930" reactiontime="+17" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="New Zealand">
              <RESULTS>
                <RESULT eventid="26" place="10" lane="7" heat="2" swimtime="00:01:26.59" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.51" />
                    <SPLIT distance="50" swimtime="00:00:21.71" />
                    <SPLIT distance="75" swimtime="00:00:31.83" />
                    <SPLIT distance="100" swimtime="00:00:43.18" />
                    <SPLIT distance="125" swimtime="00:00:53.05" />
                    <SPLIT distance="150" swimtime="00:01:04.75" />
                    <SPLIT distance="175" swimtime="00:01:15.12" />
                    <SPLIT distance="200" swimtime="00:01:26.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202034" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="202035" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="161935" reactiontime="+16" />
                    <RELAYPOSITION number="4" athleteid="214488" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="New Zealand">
              <RESULTS>
                <RESULT eventid="127" place="7" lane="7" heat="1" swimtime="00:01:30.38" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.36" />
                    <SPLIT distance="50" swimtime="00:00:21.52" />
                    <SPLIT distance="75" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:00:42.27" />
                    <SPLIT distance="125" swimtime="00:00:53.44" />
                    <SPLIT distance="150" swimtime="00:01:06.37" />
                    <SPLIT distance="175" swimtime="00:01:17.64" />
                    <SPLIT distance="200" swimtime="00:01:30.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202035" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="202034" reactiontime="+14" />
                    <RELAYPOSITION number="3" athleteid="156796" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="156788" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="6" lane="7" heat="1" swimtime="00:01:31.39" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.44" />
                    <SPLIT distance="50" swimtime="00:00:21.65" />
                    <SPLIT distance="75" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:00:42.97" />
                    <SPLIT distance="125" swimtime="00:00:54.17" />
                    <SPLIT distance="150" swimtime="00:01:06.93" />
                    <SPLIT distance="175" swimtime="00:01:18.35" />
                    <SPLIT distance="200" swimtime="00:01:31.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202035" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="161935" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="156796" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="156788" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="New Zealand">
              <RESULTS>
                <RESULT eventid="8" place="12" lane="1" heat="1" swimtime="00:03:40.47" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                    <SPLIT distance="75" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:00:54.56" />
                    <SPLIT distance="125" swimtime="00:01:06.12" />
                    <SPLIT distance="150" swimtime="00:01:19.52" />
                    <SPLIT distance="175" swimtime="00:01:33.56" />
                    <SPLIT distance="200" swimtime="00:01:47.85" />
                    <SPLIT distance="225" swimtime="00:02:00.23" />
                    <SPLIT distance="250" swimtime="00:02:14.45" />
                    <SPLIT distance="275" swimtime="00:02:29.50" />
                    <SPLIT distance="300" swimtime="00:02:44.39" />
                    <SPLIT distance="325" swimtime="00:02:56.90" />
                    <SPLIT distance="350" swimtime="00:03:11.27" />
                    <SPLIT distance="375" swimtime="00:03:26.04" />
                    <SPLIT distance="400" swimtime="00:03:40.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156788" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="156796" reactiontime="+35" />
                    <RELAYPOSITION number="3" athleteid="156844" reactiontime="+48" />
                    <RELAYPOSITION number="4" athleteid="212854" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="New Zealand">
              <RESULTS>
                <RESULT eventid="47" place="13" lane="1" heat="1" swimtime="00:04:00.92" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                    <SPLIT distance="75" swimtime="00:00:44.13" />
                    <SPLIT distance="100" swimtime="00:01:00.01" />
                    <SPLIT distance="125" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:01:31.13" />
                    <SPLIT distance="175" swimtime="00:01:48.47" />
                    <SPLIT distance="200" swimtime="00:02:06.78" />
                    <SPLIT distance="225" swimtime="00:02:18.57" />
                    <SPLIT distance="250" swimtime="00:02:33.72" />
                    <SPLIT distance="275" swimtime="00:02:49.84" />
                    <SPLIT distance="300" swimtime="00:03:06.79" />
                    <SPLIT distance="325" swimtime="00:03:18.45" />
                    <SPLIT distance="350" swimtime="00:03:32.00" />
                    <SPLIT distance="375" swimtime="00:03:46.23" />
                    <SPLIT distance="400" swimtime="00:04:00.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156788" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="143885" reactiontime="+37" />
                    <RELAYPOSITION number="3" athleteid="156844" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="156796" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="New Zealand">
              <RESULTS>
                <RESULT eventid="117" place="8" lane="8" heat="1" swimtime="00:07:50.76" reactiontime="+73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="75" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:00:55.90" />
                    <SPLIT distance="125" swimtime="00:01:10.79" />
                    <SPLIT distance="150" swimtime="00:01:25.75" />
                    <SPLIT distance="175" swimtime="00:01:40.41" />
                    <SPLIT distance="200" swimtime="00:01:54.46" />
                    <SPLIT distance="225" swimtime="00:02:06.95" />
                    <SPLIT distance="250" swimtime="00:02:21.54" />
                    <SPLIT distance="275" swimtime="00:02:36.30" />
                    <SPLIT distance="300" swimtime="00:02:51.16" />
                    <SPLIT distance="325" swimtime="00:03:06.20" />
                    <SPLIT distance="350" swimtime="00:03:21.42" />
                    <SPLIT distance="375" swimtime="00:03:36.72" />
                    <SPLIT distance="400" swimtime="00:03:51.60" />
                    <SPLIT distance="425" swimtime="00:04:04.39" />
                    <SPLIT distance="450" swimtime="00:04:19.20" />
                    <SPLIT distance="475" swimtime="00:04:34.40" />
                    <SPLIT distance="500" swimtime="00:04:49.73" />
                    <SPLIT distance="525" swimtime="00:05:05.34" />
                    <SPLIT distance="550" swimtime="00:05:20.98" />
                    <SPLIT distance="575" swimtime="00:05:36.89" />
                    <SPLIT distance="600" swimtime="00:05:52.32" />
                    <SPLIT distance="625" swimtime="00:06:05.11" />
                    <SPLIT distance="650" swimtime="00:06:19.67" />
                    <SPLIT distance="675" swimtime="00:06:34.75" />
                    <SPLIT distance="700" swimtime="00:06:50.03" />
                    <SPLIT distance="725" swimtime="00:07:05.30" />
                    <SPLIT distance="750" swimtime="00:07:20.63" />
                    <SPLIT distance="775" swimtime="00:07:35.96" />
                    <SPLIT distance="800" swimtime="00:07:50.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="161792" reactiontime="+73" />
                    <RELAYPOSITION number="2" athleteid="156786" reactiontime="+11" />
                    <RELAYPOSITION number="3" athleteid="212854" reactiontime="+14" />
                    <RELAYPOSITION number="4" athleteid="202036" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="8" lane="2" heat="2" swimtime="00:07:50.73" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.61" />
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                    <SPLIT distance="75" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:00:55.60" />
                    <SPLIT distance="125" swimtime="00:01:10.32" />
                    <SPLIT distance="150" swimtime="00:01:25.37" />
                    <SPLIT distance="175" swimtime="00:01:40.12" />
                    <SPLIT distance="200" swimtime="00:01:54.24" />
                    <SPLIT distance="225" swimtime="00:02:07.17" />
                    <SPLIT distance="250" swimtime="00:02:21.74" />
                    <SPLIT distance="275" swimtime="00:02:36.69" />
                    <SPLIT distance="300" swimtime="00:02:51.87" />
                    <SPLIT distance="325" swimtime="00:03:06.84" />
                    <SPLIT distance="350" swimtime="00:03:22.07" />
                    <SPLIT distance="375" swimtime="00:03:37.19" />
                    <SPLIT distance="400" swimtime="00:03:51.78" />
                    <SPLIT distance="425" swimtime="00:04:04.54" />
                    <SPLIT distance="450" swimtime="00:04:19.29" />
                    <SPLIT distance="475" swimtime="00:04:34.29" />
                    <SPLIT distance="500" swimtime="00:04:49.66" />
                    <SPLIT distance="525" swimtime="00:05:04.96" />
                    <SPLIT distance="550" swimtime="00:05:20.44" />
                    <SPLIT distance="575" swimtime="00:05:36.07" />
                    <SPLIT distance="600" swimtime="00:05:51.36" />
                    <SPLIT distance="625" swimtime="00:06:03.99" />
                    <SPLIT distance="650" swimtime="00:06:18.57" />
                    <SPLIT distance="675" swimtime="00:06:33.33" />
                    <SPLIT distance="700" swimtime="00:06:48.52" />
                    <SPLIT distance="725" swimtime="00:07:03.93" />
                    <SPLIT distance="750" swimtime="00:07:19.60" />
                    <SPLIT distance="775" swimtime="00:07:35.33" />
                    <SPLIT distance="800" swimtime="00:07:50.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="161792" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="156786" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="212854" reactiontime="+4" />
                    <RELAYPOSITION number="4" athleteid="202036" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="New Zealand">
              <RESULTS>
                <RESULT eventid="125" place="8" lane="8" heat="1" swimtime="00:01:37.93" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:24.82" />
                    <SPLIT distance="75" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:00:48.95" />
                    <SPLIT distance="125" swimtime="00:01:00.35" />
                    <SPLIT distance="150" swimtime="00:01:13.35" />
                    <SPLIT distance="175" swimtime="00:01:25.04" />
                    <SPLIT distance="200" swimtime="00:01:37.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="143885" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="156796" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="156788" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="161792" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="8" lane="7" heat="2" swimtime="00:01:38.45" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="75" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:00:49.09" />
                    <SPLIT distance="125" swimtime="00:01:00.45" />
                    <SPLIT distance="150" swimtime="00:01:13.47" />
                    <SPLIT distance="175" swimtime="00:01:25.41" />
                    <SPLIT distance="200" swimtime="00:01:38.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="143885" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="156796" reactiontime="+8" />
                    <RELAYPOSITION number="3" athleteid="156788" reactiontime="+17" />
                    <RELAYPOSITION number="4" athleteid="161792" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="New Zealand">
              <RESULTS>
                <RESULT eventid="11" place="11" lane="1" heat="2" swimtime="00:01:39.53" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:24.07" />
                    <SPLIT distance="75" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:00:50.18" />
                    <SPLIT distance="125" swimtime="00:01:01.56" />
                    <SPLIT distance="150" swimtime="00:01:15.57" />
                    <SPLIT distance="175" swimtime="00:01:26.75" />
                    <SPLIT distance="200" swimtime="00:01:39.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="161935" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="212856" reactiontime="+15" />
                    <RELAYPOSITION number="3" athleteid="143885" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="156796" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="New Zealand">
              <RESULTS>
                <RESULT eventid="35" place="12" lane="5" heat="1" swimtime="00:01:34.86" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.64" />
                    <SPLIT distance="50" swimtime="00:00:24.39" />
                    <SPLIT distance="75" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:00:50.87" />
                    <SPLIT distance="125" swimtime="00:01:00.97" />
                    <SPLIT distance="150" swimtime="00:01:13.43" />
                    <SPLIT distance="175" swimtime="00:01:23.53" />
                    <SPLIT distance="200" swimtime="00:01:34.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="161935" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="212856" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="202034" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="202035" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Oman" shortname="OMA" code="OMA" nation="OMA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="108528" lastname="AL ADAWI" firstname="Issa Samir Hamed" gender="M" birthdate="1999-03-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.81" eventid="14" heat="4" lane="5">
                  <MEETINFO date="2021-07-27" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.57" eventid="31" heat="4" lane="3">
                  <MEETINFO date="2021-07-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="59" lane="5" heat="4" heatid="40014" swimtime="00:00:51.05" reactiontime="+62" points="677">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                    <SPLIT distance="50" swimtime="00:00:23.98" />
                    <SPLIT distance="75" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:00:51.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="52" lane="3" heat="4" heatid="40031" swimtime="00:00:23.60" reactiontime="+66" points="623">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                    <SPLIT distance="50" swimtime="00:00:23.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Pakistan" shortname="PAK" code="PAK" nation="PAK" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="213965" lastname="KHAN" firstname="Shahbaz" gender="M" birthdate="1991-08-25">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5" heat="1" lane="5" />
                <ENTRY entrytime="NT" eventid="31" heat="2" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="60" lane="5" heat="1" heatid="10005" swimtime="00:00:27.41" reactiontime="+66" points="499">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="66" lane="8" heat="2" heatid="20031" swimtime="00:00:25.16" reactiontime="+71" points="514">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="193195" lastname="NABI" firstname="Jehanara" gender="F" birthdate="2004-07-14">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.16" eventid="43" heat="1" lane="5">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:04:28.88" eventid="1" heat="1" lane="6">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="30" lane="5" heat="1" heatid="10043" swimtime="00:02:06.32" reactiontime="+71" points="665">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                    <SPLIT distance="75" swimtime="00:00:45.23" />
                    <SPLIT distance="100" swimtime="00:01:01.36" />
                    <SPLIT distance="125" swimtime="00:01:17.46" />
                    <SPLIT distance="150" swimtime="00:01:34.00" />
                    <SPLIT distance="175" swimtime="00:01:50.52" />
                    <SPLIT distance="200" swimtime="00:02:06.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="25" lane="6" heat="1" heatid="10001" swimtime="00:04:25.36" reactiontime="+72" points="685">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="75" swimtime="00:00:45.88" />
                    <SPLIT distance="100" swimtime="00:01:02.83" />
                    <SPLIT distance="125" swimtime="00:01:19.59" />
                    <SPLIT distance="150" swimtime="00:01:36.31" />
                    <SPLIT distance="175" swimtime="00:01:52.88" />
                    <SPLIT distance="200" swimtime="00:02:09.71" />
                    <SPLIT distance="225" swimtime="00:02:26.65" />
                    <SPLIT distance="250" swimtime="00:02:43.77" />
                    <SPLIT distance="275" swimtime="00:03:00.88" />
                    <SPLIT distance="300" swimtime="00:03:18.16" />
                    <SPLIT distance="325" swimtime="00:03:35.26" />
                    <SPLIT distance="350" swimtime="00:03:52.31" />
                    <SPLIT distance="375" swimtime="00:04:09.15" />
                    <SPLIT distance="400" swimtime="00:04:25.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Panama" shortname="PAN" code="PAN" nation="PAN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="110920" lastname="CALDERON HARPER" firstname="Jeancarlo" gender="M" birthdate="1999-07-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.84" eventid="14" heat="4" lane="3">
                  <MEETINFO date="2022-10-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="44" heat="1" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="54" lane="3" heat="4" heatid="40014" swimtime="00:00:50.54" reactiontime="+58" points="698">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.36" />
                    <SPLIT distance="50" swimtime="00:00:24.37" />
                    <SPLIT distance="75" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:00:50.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="-1" lane="8" heat="1" heatid="10044" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156718" lastname="CASTILLO" firstname="Maria" gender="F" birthdate="2003-04-21">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="13" heat="2" lane="7" />
                <ENTRY entrytime="NT" eventid="4" heat="1" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="43" lane="7" heat="2" heatid="20013" swimtime="00:00:57.58" reactiontime="+73" points="664">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="75" swimtime="00:00:42.36" />
                    <SPLIT distance="100" swimtime="00:00:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="-1" lane="2" heat="1" heatid="10004" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140102" lastname="CERMELLI" firstname="Carolina" gender="F" birthdate="2001-01-31">
              <ENTRIES>
                <ENTRY entrytime="00:02:16.12" eventid="45" heat="1" lane="4">
                  <MEETINFO date="2021-10-09" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.90" eventid="18" heat="3" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="30" lane="4" heat="1" heatid="10045" swimtime="00:02:12.40" reactiontime="+59" points="724">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.19" />
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="75" swimtime="00:00:48.29" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="125" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:01:39.05" />
                    <SPLIT distance="175" swimtime="00:01:56.12" />
                    <SPLIT distance="200" swimtime="00:02:12.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="36" lane="3" heat="3" heatid="30018" swimtime="00:00:29.00" reactiontime="+60" points="661">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.40" />
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Paraguay" shortname="PAR" code="PAR" nation="PAR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="101927" lastname="HOCKIN BRUSQUETTI" firstname="Charles" gender="M" birthdate="1989-11-04">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.19" eventid="3" heat="3" lane="3">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:24.12" eventid="19" heat="3" lane="5">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="33" lane="3" heat="3" heatid="30003" swimtime="00:00:53.88" reactiontime="+59" points="721">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:25.63" />
                    <SPLIT distance="75" swimtime="00:00:39.87" />
                    <SPLIT distance="100" swimtime="00:00:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="28" lane="5" heat="3" heatid="30019" swimtime="00:00:24.29" reactiontime="+56" points="765">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.81" />
                    <SPLIT distance="50" swimtime="00:00:24.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101472" lastname="HOCKIN" firstname="Benjamin" gender="M" birthdate="1986-09-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.67" eventid="39" heat="3" lane="5">
                  <MEETINFO date="2022-10-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.35" eventid="14" heat="7" lane="3">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.50" eventid="5" heat="6" lane="1">
                  <MEETINFO date="2022-09-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.59" eventid="23" heat="2" lane="3">
                  <MEETINFO date="2022-09-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="39" lane="5" heat="3" heatid="30039" swimtime="00:00:53.87" reactiontime="+71" points="697">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.32" />
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                    <SPLIT distance="75" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:00:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="45" lane="3" heat="7" heatid="70014" swimtime="00:00:48.48" reactiontime="+71" points="791">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.12" />
                    <SPLIT distance="50" swimtime="00:00:23.34" />
                    <SPLIT distance="75" swimtime="00:00:35.89" />
                    <SPLIT distance="100" swimtime="00:00:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="40" lane="1" heat="6" heatid="60005" swimtime="00:00:23.32" reactiontime="+72" points="811">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.61" />
                    <SPLIT distance="50" swimtime="00:00:23.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="27" lane="3" heat="2" heatid="20023" swimtime="00:00:54.47" reactiontime="+72" points="740">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.92" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:00:54.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="125005" lastname="MATEOS" firstname="Matheo" gender="M" birthdate="2000-11-10">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.31" eventid="7" heat="1" lane="4">
                  <MEETINFO date="2022-04-02" />
                </ENTRY>
                <ENTRY entrytime="00:04:24.64" eventid="37" heat="1" lane="7">
                  <MEETINFO date="2022-10-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="-1" lane="4" heat="1" heatid="10007" swimtime="00:01:59.75" status="DSQ" reactiontime="+68" />
                <RESULT eventid="37" place="18" lane="7" heat="1" heatid="10037" swimtime="00:04:14.73" reactiontime="+73" points="783">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.35" />
                    <SPLIT distance="50" swimtime="00:00:27.51" />
                    <SPLIT distance="75" swimtime="00:00:43.15" />
                    <SPLIT distance="100" swimtime="00:00:59.03" />
                    <SPLIT distance="125" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:32.09" />
                    <SPLIT distance="175" swimtime="00:01:48.29" />
                    <SPLIT distance="200" swimtime="00:02:04.03" />
                    <SPLIT distance="225" swimtime="00:02:22.17" />
                    <SPLIT distance="250" swimtime="00:02:40.22" />
                    <SPLIT distance="275" swimtime="00:02:58.39" />
                    <SPLIT distance="300" swimtime="00:03:16.56" />
                    <SPLIT distance="325" swimtime="00:03:31.72" />
                    <SPLIT distance="350" swimtime="00:03:46.14" />
                    <SPLIT distance="375" swimtime="00:04:00.69" />
                    <SPLIT distance="400" swimtime="00:04:14.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110325" lastname="PRONO" firstname="Renato" gender="M" birthdate="1991-03-02">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:26.65" eventid="41" heat="7" lane="1">
                  <MEETINFO date="2021-10-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="24" lane="1" heat="7" heatid="70041" swimtime="00:00:26.92" reactiontime="+60" points="796">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.16" />
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130276" lastname="ALONSO" firstname="Luana" gender="F" birthdate="2004-03-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.90" eventid="38" heat="4" lane="8">
                  <MEETINFO date="2022-08-10" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.46" eventid="20" heat="3" lane="1">
                  <MEETINFO date="2022-09-15" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="22" lane="8" heat="4" heatid="40038" swimtime="00:00:58.93" reactiontime="+66" points="794">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.32" />
                    <SPLIT distance="50" swimtime="00:00:27.10" />
                    <SPLIT distance="75" swimtime="00:00:42.54" />
                    <SPLIT distance="100" swimtime="00:00:58.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="20" lane="1" heat="3" heatid="30020" swimtime="00:02:12.19" reactiontime="+69" points="740">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                    <SPLIT distance="75" swimtime="00:00:45.10" />
                    <SPLIT distance="100" swimtime="00:01:01.92" />
                    <SPLIT distance="125" swimtime="00:01:18.50" />
                    <SPLIT distance="150" swimtime="00:01:35.87" />
                    <SPLIT distance="175" swimtime="00:01:53.81" />
                    <SPLIT distance="200" swimtime="00:02:12.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Paraguay">
              <RESULTS>
                <RESULT eventid="26" place="14" lane="7" heat="1" swimtime="00:01:31.17" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.82" />
                    <SPLIT distance="50" swimtime="00:00:22.36" />
                    <SPLIT distance="75" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:00:45.39" />
                    <SPLIT distance="125" swimtime="00:00:56.52" />
                    <SPLIT distance="150" swimtime="00:01:08.63" />
                    <SPLIT distance="175" swimtime="00:01:19.16" />
                    <SPLIT distance="200" swimtime="00:01:31.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101472" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="110325" reactiontime="+48" />
                    <RELAYPOSITION number="3" athleteid="125005" reactiontime="+48" />
                    <RELAYPOSITION number="4" athleteid="101927" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Paraguay">
              <RESULTS>
                <RESULT eventid="35" place="15" lane="7" heat="2" swimtime="00:01:37.18" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:24.50" />
                    <SPLIT distance="75" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:00:51.02" />
                    <SPLIT distance="125" swimtime="00:01:01.56" />
                    <SPLIT distance="150" swimtime="00:01:14.25" />
                    <SPLIT distance="175" swimtime="00:01:25.13" />
                    <SPLIT distance="200" swimtime="00:01:37.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="101927" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="110325" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="101472" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="125005" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Peru" shortname="PER" code="PER" nation="PER" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="154229" lastname="NICOLAS MATTA" firstname="Javier Borja" gender="M" birthdate="2000-09-23">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.30" eventid="39" heat="4" lane="6">
                  <MEETINFO date="2022-10-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="23" heat="1" lane="2" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="28" lane="6" heat="4" heatid="40039" swimtime="00:00:51.77" reactiontime="+56" points="786">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.89" />
                    <SPLIT distance="50" swimtime="00:00:23.73" />
                    <SPLIT distance="75" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:00:51.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="23" lane="2" heat="1" heatid="10023" swimtime="00:00:53.75" reactiontime="+54" points="770">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:24.10" />
                    <SPLIT distance="75" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:00:53.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145014" lastname="VARGAS" firstname="Joaquin" gender="M" birthdate="2002-02-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.68" eventid="44" heat="3" lane="5">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:03:43.32" eventid="24" heat="3" lane="3">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="27" lane="5" heat="3" heatid="30044" swimtime="00:01:45.69" reactiontime="+66" points="831">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.78" />
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                    <SPLIT distance="75" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:00:51.32" />
                    <SPLIT distance="125" swimtime="00:01:04.95" />
                    <SPLIT distance="150" swimtime="00:01:18.50" />
                    <SPLIT distance="175" swimtime="00:01:32.19" />
                    <SPLIT distance="200" swimtime="00:01:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="18" lane="3" heat="3" heatid="30024" swimtime="00:03:45.66" reactiontime="+67" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.10" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:00:53.89" />
                    <SPLIT distance="125" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:22.45" />
                    <SPLIT distance="175" swimtime="00:01:36.77" />
                    <SPLIT distance="200" swimtime="00:01:51.21" />
                    <SPLIT distance="225" swimtime="00:02:05.67" />
                    <SPLIT distance="250" swimtime="00:02:19.89" />
                    <SPLIT distance="275" swimtime="00:02:34.25" />
                    <SPLIT distance="300" swimtime="00:02:48.59" />
                    <SPLIT distance="325" swimtime="00:03:02.84" />
                    <SPLIT distance="350" swimtime="00:03:17.29" />
                    <SPLIT distance="375" swimtime="00:03:31.68" />
                    <SPLIT distance="400" swimtime="00:03:45.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202805" lastname="FERNANDINI ERAZO" firstname="Rafaela" gender="F" birthdate="2001-06-17">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:55.12" eventid="13" heat="6" lane="7">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.36" eventid="30" heat="5" lane="6">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="37" lane="7" heat="6" heatid="60013" swimtime="00:00:55.70" reactiontime="+66" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.44" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                    <SPLIT distance="75" swimtime="00:00:41.12" />
                    <SPLIT distance="100" swimtime="00:00:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="29" lane="6" heat="5" heatid="50030" swimtime="00:00:25.36" reactiontime="+63" points="739">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.25" />
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196772" lastname="SOTOMAYOR" firstname="Alexia" gender="F" birthdate="2006-07-18">
              <ENTRIES>
                <ENTRY entrytime="00:02:13.80" eventid="45" heat="2" lane="7">
                  <MEETINFO date="2022-10-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:28.11" eventid="18" heat="4" lane="3">
                  <MEETINFO date="2021-10-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="29" lane="7" heat="2" heatid="20045" swimtime="00:02:12.36" reactiontime="+54" points="725">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="75" swimtime="00:00:46.81" />
                    <SPLIT distance="100" swimtime="00:01:03.67" />
                    <SPLIT distance="125" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:01:37.38" />
                    <SPLIT distance="175" swimtime="00:01:54.86" />
                    <SPLIT distance="200" swimtime="00:02:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="29" lane="3" heat="4" heatid="40018" swimtime="00:00:28.06" reactiontime="+52" points="730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="163914" lastname="MUÑOZ" firstname="Maria Fe" gender="F" birthdate="1999-06-20">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.01" eventid="20" heat="2" lane="7">
                  <MEETINFO date="2021-10-31" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="23" lane="7" heat="2" heatid="20020" swimtime="00:02:16.82" reactiontime="+69" points="668">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="75" swimtime="00:00:46.97" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="125" swimtime="00:01:21.27" />
                    <SPLIT distance="150" swimtime="00:01:39.03" />
                    <SPLIT distance="175" swimtime="00:01:57.68" />
                    <SPLIT distance="200" swimtime="00:02:16.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144565" lastname="DE BEVER" firstname="Mckenna" gender="F" birthdate="1996-06-05">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:02:11.45" eventid="6" heat="3" lane="8">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:01:00.65" eventid="22" heat="3" lane="7">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="26" lane="8" heat="3" heatid="30006" swimtime="00:02:12.85" reactiontime="+68" points="771">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="75" swimtime="00:00:45.85" />
                    <SPLIT distance="100" swimtime="00:01:02.42" />
                    <SPLIT distance="125" swimtime="00:01:21.35" />
                    <SPLIT distance="150" swimtime="00:01:40.81" />
                    <SPLIT distance="175" swimtime="00:01:57.30" />
                    <SPLIT distance="200" swimtime="00:02:12.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="17" lane="7" heat="3" heatid="30022" swimtime="00:01:00.48" reactiontime="+66" points="815">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.75" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="75" swimtime="00:00:45.74" />
                    <SPLIT distance="100" swimtime="00:01:00.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Peru">
              <RESULTS>
                <RESULT eventid="27" place="15" lane="1" heat="2" swimtime="00:01:35.41" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.50" />
                    <SPLIT distance="50" swimtime="00:00:22.05" />
                    <SPLIT distance="75" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:00:44.96" />
                    <SPLIT distance="125" swimtime="00:00:56.85" />
                    <SPLIT distance="150" swimtime="00:01:09.95" />
                    <SPLIT distance="175" swimtime="00:01:21.92" />
                    <SPLIT distance="200" swimtime="00:01:35.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154229" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="145014" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="202805" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="144565" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Peru">
              <RESULTS>
                <RESULT eventid="8" place="14" lane="1" heat="2" swimtime="00:03:47.22" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.51" />
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="75" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:00:55.43" />
                    <SPLIT distance="125" swimtime="00:01:07.99" />
                    <SPLIT distance="150" swimtime="00:01:22.07" />
                    <SPLIT distance="175" swimtime="00:01:36.60" />
                    <SPLIT distance="200" swimtime="00:01:51.11" />
                    <SPLIT distance="225" swimtime="00:02:03.54" />
                    <SPLIT distance="250" swimtime="00:02:17.95" />
                    <SPLIT distance="275" swimtime="00:02:33.24" />
                    <SPLIT distance="300" swimtime="00:02:48.97" />
                    <SPLIT distance="325" swimtime="00:03:01.90" />
                    <SPLIT distance="350" swimtime="00:03:16.71" />
                    <SPLIT distance="375" swimtime="00:03:32.00" />
                    <SPLIT distance="400" swimtime="00:03:47.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202805" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="144565" reactiontime="+38" />
                    <RELAYPOSITION number="3" athleteid="196772" reactiontime="+47" />
                    <RELAYPOSITION number="4" athleteid="163914" reactiontime="+15" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Peru">
              <RESULTS>
                <RESULT eventid="47" place="15" lane="8" heat="2" swimtime="00:04:12.73" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.34" />
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="75" swimtime="00:00:45.44" />
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                    <SPLIT distance="125" swimtime="00:01:16.38" />
                    <SPLIT distance="150" swimtime="00:01:34.48" />
                    <SPLIT distance="175" swimtime="00:01:53.23" />
                    <SPLIT distance="200" swimtime="00:02:12.70" />
                    <SPLIT distance="225" swimtime="00:02:25.85" />
                    <SPLIT distance="250" swimtime="00:02:42.08" />
                    <SPLIT distance="275" swimtime="00:02:58.75" />
                    <SPLIT distance="300" swimtime="00:03:15.91" />
                    <SPLIT distance="325" swimtime="00:03:28.30" />
                    <SPLIT distance="350" swimtime="00:03:42.82" />
                    <SPLIT distance="375" swimtime="00:03:57.93" />
                    <SPLIT distance="400" swimtime="00:04:12.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196772" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="144565" reactiontime="+6" />
                    <RELAYPOSITION number="3" athleteid="163914" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="202805" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Peru">
              <RESULTS>
                <RESULT eventid="25" place="12" lane="7" heat="1" swimtime="00:01:43.84" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:25.18" />
                    <SPLIT distance="75" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:00:50.38" />
                    <SPLIT distance="125" swimtime="00:01:03.35" />
                    <SPLIT distance="150" swimtime="00:01:17.60" />
                    <SPLIT distance="175" swimtime="00:01:30.00" />
                    <SPLIT distance="200" swimtime="00:01:43.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="202805" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="144565" reactiontime="+28" />
                    <RELAYPOSITION number="3" athleteid="163914" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="196772" reactiontime="+29" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Peru">
              <RESULTS>
                <RESULT eventid="34" place="14" lane="2" heat="1" swimtime="00:01:54.18" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.85" />
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                    <SPLIT distance="75" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:01:00.85" />
                    <SPLIT distance="125" swimtime="00:01:13.70" />
                    <SPLIT distance="150" swimtime="00:01:29.06" />
                    <SPLIT distance="175" swimtime="00:01:41.08" />
                    <SPLIT distance="200" swimtime="00:01:54.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196772" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="144565" reactiontime="+17" />
                    <RELAYPOSITION number="3" athleteid="163914" reactiontime="+32" />
                    <RELAYPOSITION number="4" athleteid="202805" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Peru">
              <RESULTS>
                <RESULT eventid="11" place="21" lane="1" heat="4" swimtime="00:01:45.80" reactiontime="+52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="75" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:00:55.22" />
                    <SPLIT distance="125" swimtime="00:01:07.67" />
                    <SPLIT distance="150" swimtime="00:01:22.87" />
                    <SPLIT distance="175" swimtime="00:01:33.84" />
                    <SPLIT distance="200" swimtime="00:01:45.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196772" reactiontime="+52" />
                    <RELAYPOSITION number="2" athleteid="154229" reactiontime="+12" />
                    <RELAYPOSITION number="3" athleteid="202805" reactiontime="+53" />
                    <RELAYPOSITION number="4" athleteid="145014" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Philippines" shortname="PHI" code="PHI" nation="PHI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="157769" lastname="COOK" firstname="Jonathan Sebastian" gender="M" birthdate="2000-04-06">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.75" eventid="16" heat="3" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:02:09.40" eventid="29" heat="2" lane="4">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="44" lane="5" heat="3" heatid="30016" swimtime="00:01:00.87" reactiontime="+63" points="749">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                    <SPLIT distance="75" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:00.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="28" lane="4" heat="2" heatid="20029" swimtime="00:02:12.91" reactiontime="+64" points="738">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="75" swimtime="00:00:46.41" />
                    <SPLIT distance="100" swimtime="00:01:03.18" />
                    <SPLIT distance="125" swimtime="00:01:20.25" />
                    <SPLIT distance="150" swimtime="00:01:37.65" />
                    <SPLIT distance="175" swimtime="00:01:55.18" />
                    <SPLIT distance="200" swimtime="00:02:12.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156722" lastname="JACINTO" firstname="Jerard" gender="M" birthdate="2001-05-05">
              <ENTRIES>
                <ENTRY entrytime="00:00:24.40" eventid="19" heat="3" lane="6">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="31" lane="6" heat="3" heatid="30019" swimtime="00:00:24.36" reactiontime="+51" points="758">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:24.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157650" lastname="ISLETA" firstname="Chloe" gender="F" birthdate="1998-05-14">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.21" eventid="2" heat="3" lane="4">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.39" eventid="45" heat="3" lane="8">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.85" eventid="6" heat="2" lane="2">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.62" eventid="18" heat="5" lane="8">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:01:01.34" eventid="22" heat="4" lane="8">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="31" lane="4" heat="3" heatid="30002" swimtime="00:01:00.25" reactiontime="+54" points="756">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.93" />
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="75" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="27" lane="8" heat="3" heatid="30045" swimtime="00:02:09.17" reactiontime="+53" points="780">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="75" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:02.84" />
                    <SPLIT distance="125" swimtime="00:01:19.31" />
                    <SPLIT distance="150" swimtime="00:01:35.55" />
                    <SPLIT distance="175" swimtime="00:01:52.29" />
                    <SPLIT distance="200" swimtime="00:02:09.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="29" lane="2" heat="2" heatid="20006" swimtime="00:02:13.77" reactiontime="+67" points="755">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.01" />
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="75" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:02.31" />
                    <SPLIT distance="125" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:01:42.04" />
                    <SPLIT distance="175" swimtime="00:01:58.73" />
                    <SPLIT distance="200" swimtime="00:02:13.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="31" lane="8" heat="5" heatid="50018" swimtime="00:00:28.08" reactiontime="+56" points="728">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.89" />
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="22" lane="8" heat="4" heatid="40022" swimtime="00:01:02.11" reactiontime="+67" points="753">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.84" />
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                    <SPLIT distance="75" swimtime="00:00:47.10" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191983" lastname="DELA CRUZ" firstname="Thanya Angelyn Cacho" gender="F" birthdate="2003-02-01">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.12" eventid="15" heat="3" lane="7">
                  <MEETINFO date="2022-10-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.35" eventid="40" heat="4" lane="8">
                  <MEETINFO date="2022-10-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="33" lane="7" heat="3" heatid="30015" swimtime="00:01:07.17" reactiontime="+60" points="800">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                    <SPLIT distance="75" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="26" lane="8" heat="4" heatid="40040" swimtime="00:00:31.19" reactiontime="+61" points="767">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102642" lastname="ALKHALDI" firstname="Jasmine" gender="F" birthdate="1993-06-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.91" eventid="13" heat="4" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.62" eventid="30" heat="5" lane="7">
                  <MEETINFO date="2022-05-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="41" lane="5" heat="4" heatid="40013" swimtime="00:00:56.51" reactiontime="+67" points="703">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                    <SPLIT distance="50" swimtime="00:00:27.35" />
                    <SPLIT distance="75" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:00:56.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="32" lane="7" heat="5" heatid="50030" swimtime="00:00:25.69" reactiontime="+69" points="711">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:25.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Philippines">
              <RESULTS>
                <RESULT eventid="27" place="-1" lane="7" heat="4" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Philippines">
              <RESULTS>
                <RESULT eventid="11" place="-1" lane="4" heat="1" status="DSQ" swimtime="00:01:44.17" reactiontime="+53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:24.26" />
                    <SPLIT distance="75" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:00:51.85" />
                    <SPLIT distance="125" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:18.75" />
                    <SPLIT distance="175" swimtime="00:01:31.14" />
                    <SPLIT distance="200" swimtime="00:01:44.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156722" reactiontime="+53" />
                    <RELAYPOSITION number="2" athleteid="157769" reactiontime="+16" status="DSQ" />
                    <RELAYPOSITION number="3" athleteid="157650" reactiontime="+24" status="DSQ" />
                    <RELAYPOSITION number="4" athleteid="102642" reactiontime="+38" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Palestine" shortname="PLE" code="PLE" nation="PLE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="191977" lastname="AL BAWWAB" firstname="Yazan" gender="M" birthdate="1999-10-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.48" eventid="3" heat="2" lane="3">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.72" eventid="19" heat="2" lane="8">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="35" lane="3" heat="2" heatid="20003" swimtime="00:00:55.23" reactiontime="+64" points="670">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.93" />
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                    <SPLIT distance="75" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:00:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="-1" lane="8" heat="2" heatid="20019" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198037" lastname="ABU GHARBIEH" firstname="Mahmoud" gender="M" birthdate="2006-03-22">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="14" heat="1" lane="1" />
                <ENTRY entrytime="00:00:24.95" eventid="31" heat="4" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="66" lane="1" heat="1" heatid="10014" swimtime="00:00:52.33" reactiontime="+67" points="629">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.95" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:00:52.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="57" lane="1" heat="4" heatid="40031" swimtime="00:00:24.20" reactiontime="+63" points="578">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:24.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182628" lastname="ABU SHAMALEH" firstname="Marina" gender="F" birthdate="2005-07-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:15.20" eventid="15" heat="2" lane="6">
                  <MEETINFO date="2022-04-14" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.00" eventid="40" heat="3" lane="6">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="45" lane="6" heat="2" heatid="20015" swimtime="00:01:13.92" reactiontime="+74" points="600">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.55" />
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="75" swimtime="00:00:53.41" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="32" lane="6" heat="3" heatid="30040" swimtime="00:00:33.49" reactiontime="+73" points="620">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.64" />
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Palau" shortname="PLW" code="PLW" nation="PLW" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="101196" lastname="DINGILIUS WALLACE" firstname="Shawn" gender="M" birthdate="1994-07-26">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.93" eventid="39" heat="2" lane="1">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.35" eventid="14" heat="2" lane="1">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="54" lane="1" heat="2" heatid="20039" swimtime="00:01:05.18" reactiontime="+77" points="393">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="75" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="81" lane="1" heat="2" heatid="20014" swimtime="00:00:58.57" reactiontime="+74" points="448">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                    <SPLIT distance="75" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:00:58.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201322" lastname="SAKURAI" firstname="Travis Dui" gender="M" birthdate="2007-05-04">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5" heat="2" lane="2" />
                <ENTRY entrytime="00:00:26.57" eventid="31" heat="3" lane="6">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="61" lane="2" heat="2" heatid="20005" swimtime="00:00:28.20" reactiontime="+67" points="458">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.00" />
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="67" lane="6" heat="3" heatid="30031" swimtime="00:00:25.57" reactiontime="+63" points="490">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:25.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213981" lastname="RULUKED" firstname="Ungilreng" gender="F" birthdate="2007-06-22">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="40" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="30" heat="2" lane="8" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="41" lane="3" heat="1" heatid="10040" swimtime="00:00:41.65" reactiontime="+64" points="322">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.00" />
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="55" lane="8" heat="2" heatid="20030" swimtime="00:00:32.04" reactiontime="+66" points="366">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.23" />
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201609" lastname="MIKEL" firstname="Galyah Ngerchesiuch" gender="F" birthdate="2006-06-09">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:39.21" eventid="4" heat="2" lane="1">
                  <MEETINFO date="2022-09-01" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="41" lane="1" heat="2" heatid="20004" swimtime="00:00:36.90" reactiontime="+75" points="288">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="30" lane="5" heat="1" heatid="10022" swimtime="00:01:22.45" reactiontime="+75" points="321">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="75" swimtime="00:01:03.49" />
                    <SPLIT distance="100" swimtime="00:01:22.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Palau">
              <RESULTS>
                <RESULT eventid="27" place="27" lane="4" heat="1" swimtime="00:01:55.93" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.25" />
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="75" swimtime="00:00:47.50" />
                    <SPLIT distance="100" swimtime="00:01:03.65" />
                    <SPLIT distance="125" swimtime="00:01:15.79" />
                    <SPLIT distance="150" swimtime="00:01:29.21" />
                    <SPLIT distance="175" swimtime="00:01:41.94" />
                    <SPLIT distance="200" swimtime="00:01:55.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="213981" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="201609" reactiontime="+41" />
                    <RELAYPOSITION number="3" athleteid="201322" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="101196" reactiontime="+46" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Papua New Guinea" shortname="PNG" code="PNG" nation="PNG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="152496" lastname="TARERE" firstname="Josh" gender="M" birthdate="2000-01-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.71" eventid="14" heat="2" lane="6">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.90" eventid="31" heat="4" lane="7">
                  <MEETINFO date="2022-06-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="74" lane="6" heat="2" heatid="20014" swimtime="00:00:54.13" reactiontime="+62" points="568">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:25.82" />
                    <SPLIT distance="75" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:00:54.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="61" lane="7" heat="4" heatid="40031" swimtime="00:00:24.35" reactiontime="+64" points="567">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:24.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213547" lastname="NOKA" firstname="Nathaniel" gender="M" birthdate="2001-07-21">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.98" eventid="41" heat="2" lane="6">
                  <MEETINFO date="2022-06-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.26" eventid="5" heat="3" lane="2">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="55" lane="6" heat="2" heatid="20041" swimtime="00:00:31.62" reactiontime="+62" points="491">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.47" />
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="58" lane="2" heat="3" heatid="30005" swimtime="00:00:26.85" reactiontime="+58" points="531">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.10" />
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106844" lastname="VELE" firstname="Georgia-Leigh" gender="F" birthdate="1998-12-11">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:01.60" eventid="13" heat="3" lane="5">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.34" eventid="4" heat="2" lane="3">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="54" lane="5" heat="3" heatid="30013" swimtime="00:01:00.93" reactiontime="+76" points="560">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.07" />
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="75" swimtime="00:00:45.44" />
                    <SPLIT distance="100" swimtime="00:01:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="35" lane="3" heat="2" heatid="20004" swimtime="00:00:29.81" reactiontime="+76" points="547">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.84" />
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213545" lastname="TOKOME-GARAP" firstname="Jhnayali" gender="F" birthdate="2008-08-26">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:02:36.44" eventid="43" heat="1" lane="7">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.33" eventid="30" heat="2" lane="6">
                  <MEETINFO date="2022-06-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="35" lane="7" heat="1" heatid="10043" swimtime="00:02:24.23" reactiontime="+66" points="447">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.19" />
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="75" swimtime="00:00:49.19" />
                    <SPLIT distance="100" swimtime="00:01:07.25" />
                    <SPLIT distance="125" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:01:45.26" />
                    <SPLIT distance="175" swimtime="00:02:05.02" />
                    <SPLIT distance="200" swimtime="00:02:24.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="45" lane="6" heat="2" heatid="20030" swimtime="00:00:28.84" reactiontime="+65" points="502">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Papua New Guinea">
              <RESULTS>
                <RESULT eventid="27" place="23" lane="3" heat="1" swimtime="00:01:45.46" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:24.36" />
                    <SPLIT distance="75" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:00:49.24" />
                    <SPLIT distance="125" swimtime="00:01:02.88" />
                    <SPLIT distance="150" swimtime="00:01:17.98" />
                    <SPLIT distance="175" swimtime="00:01:31.38" />
                    <SPLIT distance="200" swimtime="00:01:45.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="152496" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="213547" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="213545" reactiontime="+2" />
                    <RELAYPOSITION number="4" athleteid="106844" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Papua New Guinea">
              <RESULTS>
                <RESULT eventid="11" place="28" lane="5" heat="1" swimtime="00:02:00.85" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.82" />
                    <SPLIT distance="50" swimtime="00:00:29.64" />
                    <SPLIT distance="75" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:01:01.34" />
                    <SPLIT distance="125" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:01:31.66" />
                    <SPLIT distance="175" swimtime="00:01:45.36" />
                    <SPLIT distance="200" swimtime="00:02:00.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="152496" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="213547" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="106844" reactiontime="+38" />
                    <RELAYPOSITION number="4" athleteid="213545" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Poland" shortname="POL" code="POL" nation="POL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="125262" lastname="STOKOWSKI" firstname="Kacper " gender="M" birthdate="1999-01-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.63" eventid="3" heat="6" lane="5">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.59" eventid="46" heat="3" lane="7">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.98" eventid="19" heat="4" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="6" lane="5" heat="1" heatid="10103" swimtime="00:00:49.74" reactiontime="+58" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.60" />
                    <SPLIT distance="50" swimtime="00:00:23.81" />
                    <SPLIT distance="75" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="5" lane="5" heat="6" heatid="60003" swimtime="00:00:50.14" reactiontime="+59" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.47" />
                    <SPLIT distance="50" swimtime="00:00:23.86" />
                    <SPLIT distance="75" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:00:50.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="2" lane="3" heat="2" heatid="20203" swimtime="00:00:49.33" reactiontime="+56" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="75" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:00:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="17" lane="7" heat="3" heatid="30046" swimtime="00:01:53.88" reactiontime="+61" points="798">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:25.66" />
                    <SPLIT distance="75" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:00:54.06" />
                    <SPLIT distance="125" swimtime="00:01:08.40" />
                    <SPLIT distance="150" swimtime="00:01:23.50" />
                    <SPLIT distance="175" swimtime="00:01:39.00" />
                    <SPLIT distance="200" swimtime="00:01:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="3" lane="3" heat="1" heatid="10119" swimtime="00:00:22.74" reactiontime="+57" points="932">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.15" />
                    <SPLIT distance="50" swimtime="00:00:22.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="1" lane="5" heat="4" heatid="40019" swimtime="00:00:22.78" reactiontime="+56" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.16" />
                    <SPLIT distance="50" swimtime="00:00:22.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="2" lane="4" heat="2" heatid="20219" swimtime="00:00:22.74" reactiontime="+57" points="932">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:22.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202181" lastname="MASIUK" firstname="Ksawery" gender="M" birthdate="2004-12-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.23" eventid="3" heat="5" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:01:46.67" eventid="44" heat="3" lane="1">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:24.44" eventid="19" heat="3" lane="2">
                  <MEETINFO date="2022-09-02" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.33" eventid="23" heat="2" lane="4">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="14" lane="7" heat="5" heatid="50003" swimtime="00:00:50.84" reactiontime="+53" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                    <SPLIT distance="75" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:00:50.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="15" lane="1" heat="1" heatid="10203" swimtime="00:00:51.01" reactiontime="+58" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.92" />
                    <SPLIT distance="50" swimtime="00:00:24.89" />
                    <SPLIT distance="75" swimtime="00:00:38.18" />
                    <SPLIT distance="100" swimtime="00:00:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="28" lane="1" heat="3" heatid="30044" swimtime="00:01:46.51" reactiontime="+67" points="812">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:24.34" />
                    <SPLIT distance="75" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:00:51.09" />
                    <SPLIT distance="125" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:19.00" />
                    <SPLIT distance="175" swimtime="00:01:33.00" />
                    <SPLIT distance="200" swimtime="00:01:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="15" lane="2" heat="3" heatid="30019" swimtime="00:00:23.35" reactiontime="+54" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:23.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="13" lane="8" heat="2" heatid="20219" swimtime="00:00:23.29" reactiontime="+54" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.39" />
                    <SPLIT distance="50" swimtime="00:00:23.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="24" lane="4" heat="2" heatid="20023" swimtime="00:00:54.05" reactiontime="+64" points="757">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.81" />
                    <SPLIT distance="50" swimtime="00:00:23.69" />
                    <SPLIT distance="75" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191675" lastname="MAJERSKI" firstname="Jakub" gender="M" birthdate="2000-08-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.65" eventid="39" heat="8" lane="3">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:01:53.02" eventid="21" heat="3" lane="7">
                  <MEETINFO date="2021-09-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.76" eventid="5" heat="9" lane="8">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="11" lane="3" heat="8" heatid="80039" swimtime="00:00:50.30" reactiontime="+67" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.75" />
                    <SPLIT distance="50" swimtime="00:00:23.40" />
                    <SPLIT distance="75" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:00:50.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="9" lane="7" heat="2" heatid="20239" swimtime="00:00:49.86" reactiontime="+67" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.10" />
                    <SPLIT distance="75" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:00:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="14" lane="7" heat="3" heatid="30021" swimtime="00:01:52.45" reactiontime="+66" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.23" />
                    <SPLIT distance="50" swimtime="00:00:24.78" />
                    <SPLIT distance="75" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:00:53.31" />
                    <SPLIT distance="125" swimtime="00:01:07.84" />
                    <SPLIT distance="150" swimtime="00:01:22.45" />
                    <SPLIT distance="175" swimtime="00:01:37.09" />
                    <SPLIT distance="200" swimtime="00:01:52.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="22" lane="8" heat="9" heatid="90005" swimtime="00:00:22.80" reactiontime="+65" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.50" />
                    <SPLIT distance="50" swimtime="00:00:22.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150124" lastname="OSTROWSKI" firstname="Karol" gender="M" birthdate="1999-09-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.94" eventid="14" heat="9" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.57" eventid="5" heat="5" lane="6">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.17" eventid="31" heat="9" lane="6">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="19" lane="7" heat="9" heatid="90014" swimtime="00:00:47.11" reactiontime="+64" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.64" />
                    <SPLIT distance="50" swimtime="00:00:22.63" />
                    <SPLIT distance="75" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="20" lane="6" heat="5" heatid="50005" swimtime="00:00:22.71" reactiontime="+65" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.36" />
                    <SPLIT distance="50" swimtime="00:00:22.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="32" lane="6" heat="9" heatid="90031" swimtime="00:00:21.54" reactiontime="+65" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.39" />
                    <SPLIT distance="50" swimtime="00:00:21.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100852" lastname="KAWECKI" firstname="Radoslaw" gender="M" birthdate="1991-08-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:48.46" eventid="46" heat="2" lane="4">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="146" place="7" lane="8" heat="1" heatid="10146" swimtime="00:01:50.33" reactiontime="+64" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:26.90" />
                    <SPLIT distance="75" swimtime="00:00:40.95" />
                    <SPLIT distance="100" swimtime="00:00:54.98" />
                    <SPLIT distance="125" swimtime="00:01:08.95" />
                    <SPLIT distance="150" swimtime="00:01:22.46" />
                    <SPLIT distance="175" swimtime="00:01:36.37" />
                    <SPLIT distance="200" swimtime="00:01:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="8" lane="4" heat="2" heatid="20046" swimtime="00:01:50.97" reactiontime="+62" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.90" />
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                    <SPLIT distance="75" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:00:54.63" />
                    <SPLIT distance="125" swimtime="00:01:08.49" />
                    <SPLIT distance="150" swimtime="00:01:22.51" />
                    <SPLIT distance="175" swimtime="00:01:36.85" />
                    <SPLIT distance="200" swimtime="00:01:50.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213056" lastname="PISKORSKA" firstname="Adela" gender="F" birthdate="2003-11-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.67" eventid="2" heat="4" lane="7">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
                <ENTRY entrytime="00:02:05.31" eventid="45" heat="3" lane="2">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.87" eventid="18" heat="7" lane="1">
                  <MEETINFO date="2022-11-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="20" lane="7" heat="4" heatid="40002" swimtime="00:00:57.74" reactiontime="+61" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="75" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:00:57.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="12" lane="2" heat="3" heatid="30045" swimtime="00:02:05.05" reactiontime="+60" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.77" />
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                    <SPLIT distance="75" swimtime="00:00:44.42" />
                    <SPLIT distance="100" swimtime="00:01:00.40" />
                    <SPLIT distance="125" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:32.22" />
                    <SPLIT distance="175" swimtime="00:01:48.65" />
                    <SPLIT distance="200" swimtime="00:02:05.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="19" lane="1" heat="7" heatid="70018" swimtime="00:00:26.77" reactiontime="+63" points="841">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.23" />
                    <SPLIT distance="50" swimtime="00:00:26.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165306" lastname="WASICK" firstname="Katarzyna" gender="F" birthdate="1992-03-22">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.44" eventid="13" heat="9" lane="5">
                  <MEETINFO date="2021-09-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.10" eventid="30" heat="8" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="8" lane="5" heat="9" heatid="90013" swimtime="00:00:52.56" reactiontime="+75" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.79" />
                    <SPLIT distance="50" swimtime="00:00:25.01" />
                    <SPLIT distance="75" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:00:52.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="9" lane="2" heat="2" heatid="20213" swimtime="00:00:52.40" reactiontime="+67" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:00:52.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="2" lane="4" heat="1" heatid="10130" swimtime="00:00:23.55" reactiontime="+68" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:23.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="1" lane="4" heat="8" heatid="80030" swimtime="00:00:23.74" reactiontime="+64" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:23.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="1" lane="4" heat="2" heatid="20230" swimtime="00:00:23.37" reactiontime="+62" points="944">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.30" />
                    <SPLIT distance="50" swimtime="00:00:23.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202173" lastname="BERNAT" firstname="Laura" gender="F" birthdate="2005-09-28">
              <ENTRIES>
                <ENTRY entrytime="00:02:05.18" eventid="45" heat="4" lane="2">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="16" lane="2" heat="4" heatid="40045" swimtime="00:02:05.54" reactiontime="+63" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.64" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:46.18" />
                    <SPLIT distance="100" swimtime="00:01:02.16" />
                    <SPLIT distance="125" swimtime="00:01:18.17" />
                    <SPLIT distance="150" swimtime="00:01:34.15" />
                    <SPLIT distance="175" swimtime="00:01:50.07" />
                    <SPLIT distance="200" swimtime="00:02:05.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Poland">
              <RESULTS>
                <RESULT eventid="26" place="-1" lane="3" heat="2" status="DSQ" swimtime="00:01:24.59" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.30" />
                    <SPLIT distance="50" swimtime="00:00:21.39" />
                    <SPLIT distance="75" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:00:42.45" />
                    <SPLIT distance="125" swimtime="00:00:52.51" />
                    <SPLIT distance="150" swimtime="00:01:03.71" />
                    <SPLIT distance="175" swimtime="00:01:13.46" />
                    <SPLIT distance="200" swimtime="00:01:24.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150124" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="191675" reactiontime="-4" status="DSQ" />
                    <RELAYPOSITION number="3" athleteid="202181" reactiontime="+19" status="DSQ" />
                    <RELAYPOSITION number="4" athleteid="125262" reactiontime="+18" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Portugal" shortname="POR" code="POR" nation="POR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="182926" lastname="COSTA" firstname="João" gender="M" birthdate="2001-08-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.87" eventid="3" heat="3" lane="1">
                  <MEETINFO date="2022-08-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:58.68" eventid="46" heat="3" lane="8">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.51" eventid="19" heat="2" lane="2">
                  <MEETINFO date="2022-03-31" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="21" lane="1" heat="3" heatid="30003" swimtime="00:00:51.34" reactiontime="+54" points="834">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:24.48" />
                    <SPLIT distance="75" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:00:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="16" lane="8" heat="3" heatid="30046" swimtime="00:01:53.54" reactiontime="+57" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.37" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="75" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:00:55.85" />
                    <SPLIT distance="125" swimtime="00:01:10.51" />
                    <SPLIT distance="150" swimtime="00:01:25.14" />
                    <SPLIT distance="175" swimtime="00:01:39.57" />
                    <SPLIT distance="200" swimtime="00:01:53.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="23" lane="2" heat="2" heatid="20019" swimtime="00:00:23.80" reactiontime="+59" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Puerto Rico" shortname="PUR" code="PUR" nation="PUR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="102228" lastname="MORALES" firstname="Yeziel" gender="M" birthdate="1996-01-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.81" eventid="3" heat="5" lane="1">
                  <MEETINFO date="2021-10-31" />
                </ENTRY>
                <ENTRY entrytime="00:01:52.16" eventid="46" heat="4" lane="1">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:01:55.71" eventid="21" heat="4" lane="1">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.06" eventid="19" heat="3" lane="4">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="30" lane="1" heat="5" heatid="50003" swimtime="00:00:52.92" reactiontime="+52" points="761">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.16" />
                    <SPLIT distance="50" swimtime="00:00:25.39" />
                    <SPLIT distance="75" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:00:52.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="19" lane="1" heat="4" heatid="40046" swimtime="00:01:53.99" reactiontime="+53" points="795">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.73" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="75" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:00:55.30" />
                    <SPLIT distance="125" swimtime="00:01:10.18" />
                    <SPLIT distance="150" swimtime="00:01:24.97" />
                    <SPLIT distance="175" swimtime="00:01:39.66" />
                    <SPLIT distance="200" swimtime="00:01:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="19" lane="1" heat="4" heatid="40021" swimtime="00:01:56.23" reactiontime="+65" points="807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:25.74" />
                    <SPLIT distance="75" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:00:55.16" />
                    <SPLIT distance="125" swimtime="00:01:10.29" />
                    <SPLIT distance="150" swimtime="00:01:25.43" />
                    <SPLIT distance="175" swimtime="00:01:40.69" />
                    <SPLIT distance="200" swimtime="00:01:56.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="-1" lane="4" heat="3" heatid="30019" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="165760" lastname="ROMANO" firstname="Kristen Elena" gender="F" birthdate="1999-09-24">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.72" eventid="6" heat="4" lane="7">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="24" lane="7" heat="4" heatid="40006" swimtime="00:02:12.07" reactiontime="+73" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="75" swimtime="00:00:45.67" />
                    <SPLIT distance="100" swimtime="00:01:01.96" />
                    <SPLIT distance="125" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:01:39.98" />
                    <SPLIT distance="175" swimtime="00:01:56.65" />
                    <SPLIT distance="200" swimtime="00:02:12.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="21" lane="4" heat="1" heatid="10022" swimtime="00:01:01.76" reactiontime="+73" points="766">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="75" swimtime="00:00:46.46" />
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214335" lastname="BROWN" firstname="Portia" gender="F" birthdate="2000-10-05">
              <ENTRIES>
                <ENTRY entrytime="00:04:40.94" eventid="36" heat="2" lane="6">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="36" place="18" lane="6" heat="2" heatid="20036" swimtime="00:04:44.68" reactiontime="+83" points="752">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.27" />
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="75" swimtime="00:00:47.64" />
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                    <SPLIT distance="125" swimtime="00:01:23.27" />
                    <SPLIT distance="150" swimtime="00:01:41.36" />
                    <SPLIT distance="175" swimtime="00:01:59.21" />
                    <SPLIT distance="200" swimtime="00:02:16.95" />
                    <SPLIT distance="225" swimtime="00:02:37.61" />
                    <SPLIT distance="250" swimtime="00:02:57.83" />
                    <SPLIT distance="275" swimtime="00:03:17.87" />
                    <SPLIT distance="300" swimtime="00:03:38.44" />
                    <SPLIT distance="325" swimtime="00:03:55.42" />
                    <SPLIT distance="350" swimtime="00:04:11.77" />
                    <SPLIT distance="375" swimtime="00:04:28.49" />
                    <SPLIT distance="400" swimtime="00:04:44.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Qatar" shortname="QAT" code="QAT" nation="QAT" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="196848" lastname="ELGHAMRY" firstname="Abdalla" gender="M" birthdate="2007-04-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.81" eventid="3" heat="2" lane="2">
                  <MEETINFO date="2021-10-27" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.19" eventid="14" heat="3" lane="7">
                  <MEETINFO date="2021-10-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="38" lane="2" heat="2" heatid="20003" swimtime="00:00:58.72" reactiontime="+68" points="557">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="75" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:00:58.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="71" lane="7" heat="3" heatid="30014" swimtime="00:00:53.57" reactiontime="+71" points="586">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:25.68" />
                    <SPLIT distance="75" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:00:53.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Romania" shortname="ROU" code="ROU" nation="ROU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="105371" lastname="GLINTA" firstname="Robert" gender="M" birthdate="1997-04-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.31" eventid="3" heat="6" lane="4">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.74" eventid="19" heat="4" lane="4">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="28" lane="4" heat="6" heatid="60003" swimtime="00:00:52.65" reactiontime="+64" points="773">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.23" />
                    <SPLIT distance="50" swimtime="00:00:25.40" />
                    <SPLIT distance="75" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:00:52.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="-1" lane="4" heat="4" heatid="40019" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196986" lastname="POPOVICI" firstname="David" gender="M" birthdate="2004-09-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.77" eventid="14" heat="9" lane="6">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:42.12" eventid="44" heat="4" lane="3">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:03:46.08" eventid="24" heat="3" lane="7">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="114" place="4" lane="2" heat="1" heatid="10114" swimtime="00:00:45.64" reactiontime="+64" points="948">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.53" />
                    <SPLIT distance="50" swimtime="00:00:22.13" />
                    <SPLIT distance="75" swimtime="00:00:33.97" />
                    <SPLIT distance="100" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="4" lane="6" heat="9" heatid="90014" swimtime="00:00:46.15" reactiontime="+64" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.72" />
                    <SPLIT distance="50" swimtime="00:00:22.44" />
                    <SPLIT distance="75" swimtime="00:00:34.41" />
                    <SPLIT distance="100" swimtime="00:00:46.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="214" place="5" lane="5" heat="1" heatid="10214" swimtime="00:00:45.91" reactiontime="+65" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.40" />
                    <SPLIT distance="75" swimtime="00:00:34.30" />
                    <SPLIT distance="100" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="144" place="2" lane="7" heat="1" heatid="10144" swimtime="00:01:40.79" reactiontime="+65" points="958">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.90" />
                    <SPLIT distance="50" swimtime="00:00:23.18" />
                    <SPLIT distance="75" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:00:49.12" />
                    <SPLIT distance="125" swimtime="00:01:02.02" />
                    <SPLIT distance="150" swimtime="00:01:15.03" />
                    <SPLIT distance="175" swimtime="00:01:28.21" />
                    <SPLIT distance="200" swimtime="00:01:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="6" lane="3" heat="4" heatid="40044" swimtime="00:01:42.31" reactiontime="+65" points="916">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:24.00" />
                    <SPLIT distance="75" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:00:50.29" />
                    <SPLIT distance="125" swimtime="00:01:03.42" />
                    <SPLIT distance="150" swimtime="00:01:16.72" />
                    <SPLIT distance="175" swimtime="00:01:30.09" />
                    <SPLIT distance="200" swimtime="00:01:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="31" lane="7" heat="3" heatid="30024" swimtime="00:03:58.48" reactiontime="+67" points="704">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:26.45" />
                    <SPLIT distance="75" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:00:56.92" />
                    <SPLIT distance="125" swimtime="00:01:12.08" />
                    <SPLIT distance="150" swimtime="00:01:27.22" />
                    <SPLIT distance="175" swimtime="00:01:42.56" />
                    <SPLIT distance="200" swimtime="00:01:57.94" />
                    <SPLIT distance="225" swimtime="00:02:13.10" />
                    <SPLIT distance="250" swimtime="00:02:28.65" />
                    <SPLIT distance="275" swimtime="00:02:43.88" />
                    <SPLIT distance="300" swimtime="00:02:58.71" />
                    <SPLIT distance="325" swimtime="00:03:13.73" />
                    <SPLIT distance="350" swimtime="00:03:29.02" />
                    <SPLIT distance="375" swimtime="00:03:44.23" />
                    <SPLIT distance="400" swimtime="00:03:58.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214216" lastname="ANGHEL" firstname="Andrei-Mircea" gender="M" birthdate="1998-07-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.14" eventid="19" heat="3" lane="8">
                  <MEETINFO date="2022-08-14" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="5" heat="2" lane="6" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="7" lane="8" heat="3" heatid="30019" swimtime="00:00:23.12" reactiontime="+55" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="-1" lane="6" heat="2" heatid="20219" swimtime="00:00:23.24" status="DSQ" reactiontime="+58" />
                <RESULT eventid="5" place="49" lane="6" heat="2" heatid="20005" swimtime="00:00:23.85" reactiontime="+62" points="758">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.73" />
                    <SPLIT distance="50" swimtime="00:00:23.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="South Africa" shortname="RSA" code="RSA" nation="RSA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="170357" lastname="COETZE" firstname="Pieter" gender="M" birthdate="2004-05-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.86" eventid="3" heat="6" lane="2">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.36" eventid="46" heat="2" lane="2">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.13" eventid="19" heat="5" lane="3">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.99" eventid="31" heat="7" lane="7">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="4" lane="7" heat="1" heatid="10103" swimtime="00:00:49.60" reactiontime="+62" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.45" />
                    <SPLIT distance="50" swimtime="00:00:24.07" />
                    <SPLIT distance="75" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:00:49.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="9" lane="2" heat="6" heatid="60003" swimtime="00:00:50.26" reactiontime="+63" points="889">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.18" />
                    <SPLIT distance="75" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:00:50.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="6" lane="2" heat="2" heatid="20203" swimtime="00:00:49.85" reactiontime="+64" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:24.00" />
                    <SPLIT distance="75" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:00:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="10" lane="2" heat="2" heatid="20046" swimtime="00:01:51.51" reactiontime="+67" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                    <SPLIT distance="75" swimtime="00:00:40.58" />
                    <SPLIT distance="100" swimtime="00:00:55.07" />
                    <SPLIT distance="125" swimtime="00:01:09.37" />
                    <SPLIT distance="150" swimtime="00:01:23.85" />
                    <SPLIT distance="175" swimtime="00:01:37.95" />
                    <SPLIT distance="200" swimtime="00:01:51.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="5" lane="6" heat="1" heatid="10119" swimtime="00:00:22.84" reactiontime="+64" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="3" lane="3" heat="5" heatid="50019" swimtime="00:00:23.01" reactiontime="+65" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:23.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="4" lane="5" heat="2" heatid="20219" swimtime="00:00:22.86" reactiontime="+64" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.28" />
                    <SPLIT distance="50" swimtime="00:00:22.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="40" lane="7" heat="7" heatid="70031" swimtime="00:00:21.68" reactiontime="+69" points="804">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.55" />
                    <SPLIT distance="50" swimtime="00:00:21.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197938" lastname="KEYLOCK" firstname="Kian" gender="M" birthdate="2005-06-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.98" eventid="16" heat="3" lane="6">
                  <MEETINFO date="2021-09-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.65" eventid="29" heat="2" lane="2">
                  <MEETINFO date="2021-09-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="43" lane="6" heat="3" heatid="30016" swimtime="00:01:00.60" reactiontime="+64" points="759">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="75" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:00.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="24" lane="2" heat="2" heatid="20029" swimtime="00:02:11.20" reactiontime="+64" points="768">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.98" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:46.91" />
                    <SPLIT distance="100" swimtime="00:01:03.40" />
                    <SPLIT distance="125" swimtime="00:01:20.04" />
                    <SPLIT distance="150" swimtime="00:01:36.83" />
                    <SPLIT distance="175" swimtime="00:01:54.00" />
                    <SPLIT distance="200" swimtime="00:02:11.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102602" lastname="LE CLOS" firstname="Chad" gender="M" birthdate="1992-04-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.58" eventid="39" heat="8" lane="4">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:49.62" eventid="21" heat="4" lane="5">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.21" eventid="5" heat="8" lane="5">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="1" lane="4" heat="1" heatid="10139" swimtime="00:00:48.59" reactiontime="+60" points="950">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.28" />
                    <SPLIT distance="50" swimtime="00:00:22.50" />
                    <SPLIT distance="75" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:00:48.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="6" lane="4" heat="8" heatid="80039" swimtime="00:00:49.88" reactiontime="+84" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.81" />
                    <SPLIT distance="50" swimtime="00:00:23.19" />
                    <SPLIT distance="75" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:00:49.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="1" lane="3" heat="1" heatid="10239" swimtime="00:00:48.98" reactiontime="+62" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.37" />
                    <SPLIT distance="50" swimtime="00:00:22.66" />
                    <SPLIT distance="75" swimtime="00:00:35.47" />
                    <SPLIT distance="100" swimtime="00:00:48.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="121" place="1" lane="5" heat="1" heatid="10121" swimtime="00:01:48.27" reactiontime="+62" points="999">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.95" />
                    <SPLIT distance="50" swimtime="00:00:24.42" />
                    <SPLIT distance="75" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:00:52.39" />
                    <SPLIT distance="125" swimtime="00:01:06.48" />
                    <SPLIT distance="150" swimtime="00:01:20.49" />
                    <SPLIT distance="175" swimtime="00:01:34.45" />
                    <SPLIT distance="200" swimtime="00:01:48.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="2" lane="5" heat="4" heatid="40021" swimtime="00:01:49.98" reactiontime="+64" points="953">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.11" />
                    <SPLIT distance="50" swimtime="00:00:24.77" />
                    <SPLIT distance="75" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:00:53.10" />
                    <SPLIT distance="125" swimtime="00:01:07.69" />
                    <SPLIT distance="150" swimtime="00:01:21.81" />
                    <SPLIT distance="175" swimtime="00:01:35.88" />
                    <SPLIT distance="200" swimtime="00:01:49.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="105" place="5" lane="2" heat="1" heatid="10105" swimtime="00:00:22.11" reactiontime="+60" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.18" />
                    <SPLIT distance="50" swimtime="00:00:22.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="7" lane="5" heat="8" heatid="80005" swimtime="00:00:22.31" reactiontime="+59" points="926">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.26" />
                    <SPLIT distance="50" swimtime="00:00:22.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="5" lane="6" heat="2" heatid="20205" swimtime="00:00:22.09" reactiontime="+61" points="954">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:22.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108867" lastname="JIMMIE" firstname="Clayton" gender="M" birthdate="1995-07-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.31" eventid="14" heat="7" lane="5">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.54" eventid="5" heat="5" lane="5">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="40" lane="5" heat="7" heatid="70014" swimtime="00:00:48.09" reactiontime="+72" points="810">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.19" />
                    <SPLIT distance="50" swimtime="00:00:23.26" />
                    <SPLIT distance="75" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:00:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="43" lane="5" heat="5" heatid="50005" swimtime="00:00:23.41" reactiontime="+69" points="801">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.59" />
                    <SPLIT distance="50" swimtime="00:00:23.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154863" lastname="SATES" firstname="Matthew" gender="M" birthdate="2003-07-28">
              <ENTRIES>
                <ENTRY entrytime="00:01:40.65" eventid="44" heat="6" lane="4">
                  <MEETINFO date="2021-10-03" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.45" eventid="7" heat="4" lane="5">
                  <MEETINFO date="2021-10-02" />
                </ENTRY>
                <ENTRY entrytime="00:03:36.30" eventid="24" heat="5" lane="5">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:04:01.98" eventid="37" heat="3" lane="6">
                  <MEETINFO date="2021-10-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="13" lane="4" heat="6" heatid="60044" swimtime="00:01:43.22" reactiontime="+66" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.31" />
                    <SPLIT distance="50" swimtime="00:00:24.22" />
                    <SPLIT distance="75" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:00:50.68" />
                    <SPLIT distance="125" swimtime="00:01:03.82" />
                    <SPLIT distance="150" swimtime="00:01:16.99" />
                    <SPLIT distance="175" swimtime="00:01:30.33" />
                    <SPLIT distance="200" swimtime="00:01:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="107" place="1" lane="6" heat="1" heatid="10107" swimtime="00:01:50.15" reactiontime="+65" points="985">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.70" />
                    <SPLIT distance="50" swimtime="00:00:23.56" />
                    <SPLIT distance="75" swimtime="00:00:37.92" />
                    <SPLIT distance="100" swimtime="00:00:51.53" />
                    <SPLIT distance="125" swimtime="00:01:07.25" />
                    <SPLIT distance="150" swimtime="00:01:23.23" />
                    <SPLIT distance="175" swimtime="00:01:37.17" />
                    <SPLIT distance="200" swimtime="00:01:50.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="4" lane="5" heat="4" heatid="40007" swimtime="00:01:52.52" reactiontime="+67" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.66" />
                    <SPLIT distance="50" swimtime="00:00:23.64" />
                    <SPLIT distance="75" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:00:52.43" />
                    <SPLIT distance="125" swimtime="00:01:08.81" />
                    <SPLIT distance="150" swimtime="00:01:25.21" />
                    <SPLIT distance="175" swimtime="00:01:39.40" />
                    <SPLIT distance="200" swimtime="00:01:52.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="12" lane="5" heat="5" heatid="50024" swimtime="00:03:41.05" reactiontime="+67" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:24.83" />
                    <SPLIT distance="75" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:00:52.32" />
                    <SPLIT distance="125" swimtime="00:01:06.03" />
                    <SPLIT distance="150" swimtime="00:01:19.78" />
                    <SPLIT distance="175" swimtime="00:01:33.78" />
                    <SPLIT distance="200" swimtime="00:01:47.72" />
                    <SPLIT distance="225" swimtime="00:02:01.74" />
                    <SPLIT distance="250" swimtime="00:02:15.52" />
                    <SPLIT distance="275" swimtime="00:02:29.24" />
                    <SPLIT distance="300" swimtime="00:02:43.23" />
                    <SPLIT distance="325" swimtime="00:02:57.26" />
                    <SPLIT distance="350" swimtime="00:03:11.57" />
                    <SPLIT distance="375" swimtime="00:03:26.49" />
                    <SPLIT distance="400" swimtime="00:03:41.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="3" lane="3" heat="1" heatid="10137" swimtime="00:03:59.21" reactiontime="+68" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.09" />
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                    <SPLIT distance="75" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:00:53.40" />
                    <SPLIT distance="125" swimtime="00:01:09.13" />
                    <SPLIT distance="150" swimtime="00:01:24.41" />
                    <SPLIT distance="175" swimtime="00:01:39.74" />
                    <SPLIT distance="200" swimtime="00:01:55.30" />
                    <SPLIT distance="225" swimtime="00:02:11.86" />
                    <SPLIT distance="250" swimtime="00:02:28.52" />
                    <SPLIT distance="275" swimtime="00:02:45.47" />
                    <SPLIT distance="300" swimtime="00:03:02.95" />
                    <SPLIT distance="325" swimtime="00:03:17.50" />
                    <SPLIT distance="350" swimtime="00:03:31.47" />
                    <SPLIT distance="375" swimtime="00:03:45.57" />
                    <SPLIT distance="400" swimtime="00:03:59.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="3" lane="6" heat="3" heatid="30037" swimtime="00:04:02.18" reactiontime="+68" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.22" />
                    <SPLIT distance="50" swimtime="00:00:24.89" />
                    <SPLIT distance="75" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:00:54.08" />
                    <SPLIT distance="125" swimtime="00:01:10.08" />
                    <SPLIT distance="150" swimtime="00:01:25.39" />
                    <SPLIT distance="175" swimtime="00:01:40.99" />
                    <SPLIT distance="200" swimtime="00:01:56.47" />
                    <SPLIT distance="225" swimtime="00:02:13.66" />
                    <SPLIT distance="250" swimtime="00:02:30.84" />
                    <SPLIT distance="275" swimtime="00:02:47.92" />
                    <SPLIT distance="300" swimtime="00:03:05.44" />
                    <SPLIT distance="325" swimtime="00:03:20.51" />
                    <SPLIT distance="350" swimtime="00:03:34.71" />
                    <SPLIT distance="375" swimtime="00:03:48.89" />
                    <SPLIT distance="400" swimtime="00:04:02.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="212656" lastname="HADDON" firstname="Simon" gender="M" birthdate="1998-10-01">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:27.74" eventid="41" heat="5" lane="8">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:54.82" eventid="23" heat="2" lane="2">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="38" lane="8" heat="5" heatid="50041" swimtime="00:00:27.67" reactiontime="+76" points="733">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.55" />
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="29" lane="2" heat="2" heatid="20023" swimtime="00:00:54.79" reactiontime="+68" points="727">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.00" />
                    <SPLIT distance="50" swimtime="00:00:24.95" />
                    <SPLIT distance="75" swimtime="00:00:41.13" />
                    <SPLIT distance="100" swimtime="00:00:54.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="210937" lastname="DRAKOPOULOS" firstname="Milla" gender="F" birthdate="2006-07-03">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:00.03" eventid="2" heat="3" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:29.00" eventid="18" heat="4" lane="1">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="36" lane="7" heat="3" heatid="30002" swimtime="00:01:01.52" reactiontime="+66" points="710">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.28" />
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="75" swimtime="00:00:45.60" />
                    <SPLIT distance="100" swimtime="00:01:01.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="31" lane="1" heat="4" heatid="40018" swimtime="00:00:28.08" reactiontime="+67" points="728">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170587" lastname="VAN NIEKERK" firstname="Lara" gender="F" birthdate="2003-05-13">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.89" eventid="15" heat="5" lane="6">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.62" eventid="40" heat="6" lane="3">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="5" lane="2" heat="1" heatid="10115" swimtime="00:01:04.12" reactiontime="+71" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.71" />
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="75" swimtime="00:00:46.65" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="2" lane="6" heat="5" heatid="50015" swimtime="00:01:03.93" reactiontime="+73" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="75" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="5" lane="4" heat="1" heatid="10215" swimtime="00:01:04.36" reactiontime="+70" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="75" swimtime="00:00:46.90" />
                    <SPLIT distance="100" swimtime="00:01:04.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="2" lane="3" heat="1" heatid="10140" swimtime="00:00:29.09" reactiontime="+68" points="946">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="3" lane="3" heat="6" heatid="60040" swimtime="00:00:29.45" reactiontime="+69" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="3" lane="5" heat="2" heatid="20240" swimtime="00:00:29.27" reactiontime="+72" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="144092" lastname="MEDER" firstname="Rebecca" gender="F" birthdate="2002-07-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.93" eventid="38" heat="4" lane="1">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.37" eventid="28" heat="3" lane="8">
                  <MEETINFO date="2022-08-14" />
                </ENTRY>
                <ENTRY entrytime="00:02:12.01" eventid="6" heat="2" lane="5">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:01:00.00" eventid="22" heat="2" lane="6">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="19" lane="1" heat="4" heatid="40038" swimtime="00:00:58.04" reactiontime="+73" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.08" />
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                    <SPLIT distance="75" swimtime="00:00:42.19" />
                    <SPLIT distance="100" swimtime="00:00:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="19" lane="8" heat="3" heatid="30028" swimtime="00:02:23.64" reactiontime="+77" points="822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="75" swimtime="00:00:51.19" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="125" swimtime="00:01:27.86" />
                    <SPLIT distance="150" swimtime="00:01:46.58" />
                    <SPLIT distance="175" swimtime="00:02:05.02" />
                    <SPLIT distance="200" swimtime="00:02:23.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="10" lane="5" heat="2" heatid="20006" swimtime="00:02:07.47" reactiontime="+72" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:27.30" />
                    <SPLIT distance="75" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:00:59.33" />
                    <SPLIT distance="125" swimtime="00:01:17.54" />
                    <SPLIT distance="150" swimtime="00:01:36.33" />
                    <SPLIT distance="175" swimtime="00:01:52.50" />
                    <SPLIT distance="200" swimtime="00:02:07.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="6" lane="2" heat="1" heatid="10122" swimtime="00:00:58.46" reactiontime="+71" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:26.70" />
                    <SPLIT distance="75" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:00:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="8" lane="6" heat="2" heatid="20022" swimtime="00:00:59.38" reactiontime="+76" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.24" />
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                    <SPLIT distance="75" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:00:59.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="5" lane="6" heat="1" heatid="10222" swimtime="00:00:58.98" reactiontime="+74" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.15" />
                    <SPLIT distance="50" swimtime="00:00:27.07" />
                    <SPLIT distance="75" swimtime="00:00:44.37" />
                    <SPLIT distance="100" swimtime="00:00:58.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="191644" lastname="DE LANGE" firstname="Caitlin" gender="F" birthdate="2004-03-04">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:55.47" eventid="13" heat="5" lane="6">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.17" eventid="30" heat="5" lane="4">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="28" lane="6" heat="5" heatid="50013" swimtime="00:00:54.47" reactiontime="+67" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.30" />
                    <SPLIT distance="50" swimtime="00:00:25.92" />
                    <SPLIT distance="75" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:00:54.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="16" lane="4" heat="5" heatid="50030" swimtime="00:00:24.67" reactiontime="+63" points="802">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:24.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="15" lane="8" heat="1" heatid="10230" swimtime="00:00:24.53" reactiontime="+67" points="816">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:24.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170443" lastname="PEARSE" firstname="Hannah" gender="F" birthdate="2003-03-30">
              <ENTRIES>
                <ENTRY entrytime="00:02:09.47" eventid="45" heat="2" lane="5">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="26" lane="5" heat="2" heatid="20045" swimtime="00:02:08.84" reactiontime="+61" points="786">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.17" />
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                    <SPLIT distance="75" swimtime="00:00:47.05" />
                    <SPLIT distance="100" swimtime="00:01:03.03" />
                    <SPLIT distance="125" swimtime="00:01:19.26" />
                    <SPLIT distance="150" swimtime="00:01:35.67" />
                    <SPLIT distance="175" swimtime="00:01:52.43" />
                    <SPLIT distance="200" swimtime="00:02:08.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="108899" lastname="VISAGIE" firstname="Emily" gender="F" birthdate="1998-01-08">
              <ENTRIES>
                <ENTRY entrytime="00:02:23.20" eventid="28" heat="5" lane="8">
                  <MEETINFO date="2021-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:29.00" eventid="4" heat="3" lane="8">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="-1" lane="8" heat="5" heatid="50028" swimtime="00:02:22.92" status="DSQ" reactiontime="+72" />
                <RESULT eventid="4" place="32" lane="8" heat="3" heatid="30004" swimtime="00:00:28.39" reactiontime="+73" points="633">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197620" lastname="TUCKER" firstname="Dakota" gender="F" birthdate="2004-10-26">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.55" eventid="20" heat="2" lane="1">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
                <ENTRY entrytime="00:04:38.16" eventid="36" heat="2" lane="4">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="17" lane="1" heat="2" heatid="20020" swimtime="00:02:11.34" reactiontime="+71" points="755">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.32" />
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="75" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:02.77" />
                    <SPLIT distance="125" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:01:36.51" />
                    <SPLIT distance="175" swimtime="00:01:53.80" />
                    <SPLIT distance="200" swimtime="00:02:11.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="14" lane="4" heat="2" heatid="20036" swimtime="00:04:40.01" reactiontime="+78" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="75" swimtime="00:00:46.33" />
                    <SPLIT distance="100" swimtime="00:01:03.12" />
                    <SPLIT distance="125" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:01:37.93" />
                    <SPLIT distance="175" swimtime="00:01:55.14" />
                    <SPLIT distance="200" swimtime="00:02:12.67" />
                    <SPLIT distance="225" swimtime="00:02:32.84" />
                    <SPLIT distance="250" swimtime="00:02:52.91" />
                    <SPLIT distance="275" swimtime="00:03:13.20" />
                    <SPLIT distance="300" swimtime="00:03:33.62" />
                    <SPLIT distance="325" swimtime="00:03:50.61" />
                    <SPLIT distance="350" swimtime="00:04:07.20" />
                    <SPLIT distance="375" swimtime="00:04:23.96" />
                    <SPLIT distance="400" swimtime="00:04:40.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="195476" lastname="HOUTMAN" firstname="Stephanie" gender="F" birthdate="2002-09-30">
              <ENTRIES>
                <ENTRY entrytime="00:04:14.19" eventid="1" heat="1" lane="4">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
                <ENTRY entrytime="00:08:39.45" eventid="12" heat="1" lane="5">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="00:16:42.10" eventid="33" heat="2" lane="7">
                  <MEETINFO date="2022-08-14" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="1" place="19" lane="4" heat="1" heatid="10001" swimtime="00:04:13.16" reactiontime="+79" points="788">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.01" />
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="75" swimtime="00:00:45.02" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="125" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:01:32.60" />
                    <SPLIT distance="175" swimtime="00:01:48.66" />
                    <SPLIT distance="200" swimtime="00:02:04.72" />
                    <SPLIT distance="225" swimtime="00:02:20.49" />
                    <SPLIT distance="250" swimtime="00:02:36.56" />
                    <SPLIT distance="275" swimtime="00:02:52.69" />
                    <SPLIT distance="300" swimtime="00:03:09.11" />
                    <SPLIT distance="325" swimtime="00:03:25.44" />
                    <SPLIT distance="350" swimtime="00:03:41.86" />
                    <SPLIT distance="375" swimtime="00:03:57.72" />
                    <SPLIT distance="400" swimtime="00:04:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="15" lane="5" heat="1" heatid="10012" swimtime="00:08:39.15" reactiontime="+79" points="787">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                    <SPLIT distance="75" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:03.25" />
                    <SPLIT distance="125" swimtime="00:01:19.62" />
                    <SPLIT distance="150" swimtime="00:01:36.20" />
                    <SPLIT distance="175" swimtime="00:01:52.55" />
                    <SPLIT distance="200" swimtime="00:02:09.19" />
                    <SPLIT distance="225" swimtime="00:02:25.32" />
                    <SPLIT distance="250" swimtime="00:02:41.59" />
                    <SPLIT distance="275" swimtime="00:02:57.70" />
                    <SPLIT distance="300" swimtime="00:03:14.01" />
                    <SPLIT distance="325" swimtime="00:03:30.06" />
                    <SPLIT distance="350" swimtime="00:03:46.46" />
                    <SPLIT distance="375" swimtime="00:04:02.63" />
                    <SPLIT distance="400" swimtime="00:04:18.99" />
                    <SPLIT distance="425" swimtime="00:04:35.01" />
                    <SPLIT distance="450" swimtime="00:04:51.43" />
                    <SPLIT distance="475" swimtime="00:05:07.67" />
                    <SPLIT distance="500" swimtime="00:05:24.36" />
                    <SPLIT distance="525" swimtime="00:05:40.51" />
                    <SPLIT distance="550" swimtime="00:05:57.28" />
                    <SPLIT distance="575" swimtime="00:06:13.46" />
                    <SPLIT distance="600" swimtime="00:06:30.26" />
                    <SPLIT distance="625" swimtime="00:06:46.50" />
                    <SPLIT distance="650" swimtime="00:07:03.06" />
                    <SPLIT distance="675" swimtime="00:07:19.51" />
                    <SPLIT distance="700" swimtime="00:07:35.92" />
                    <SPLIT distance="725" swimtime="00:07:52.05" />
                    <SPLIT distance="750" swimtime="00:08:08.58" />
                    <SPLIT distance="775" swimtime="00:08:24.27" />
                    <SPLIT distance="800" swimtime="00:08:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="13" lane="7" heat="2" heatid="20033" swimtime="00:16:35.55" reactiontime="+78" points="784">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                    <SPLIT distance="75" swimtime="00:00:47.10" />
                    <SPLIT distance="100" swimtime="00:01:03.85" />
                    <SPLIT distance="125" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:01:37.33" />
                    <SPLIT distance="175" swimtime="00:01:53.93" />
                    <SPLIT distance="200" swimtime="00:02:10.71" />
                    <SPLIT distance="225" swimtime="00:02:27.23" />
                    <SPLIT distance="250" swimtime="00:02:43.95" />
                    <SPLIT distance="275" swimtime="00:03:00.53" />
                    <SPLIT distance="300" swimtime="00:03:17.31" />
                    <SPLIT distance="325" swimtime="00:03:33.88" />
                    <SPLIT distance="350" swimtime="00:03:50.63" />
                    <SPLIT distance="375" swimtime="00:04:07.13" />
                    <SPLIT distance="400" swimtime="00:04:23.74" />
                    <SPLIT distance="425" swimtime="00:04:40.25" />
                    <SPLIT distance="450" swimtime="00:04:56.99" />
                    <SPLIT distance="475" swimtime="00:05:13.23" />
                    <SPLIT distance="500" swimtime="00:05:29.67" />
                    <SPLIT distance="525" swimtime="00:05:46.08" />
                    <SPLIT distance="550" swimtime="00:06:02.86" />
                    <SPLIT distance="575" swimtime="00:06:19.25" />
                    <SPLIT distance="600" swimtime="00:06:36.06" />
                    <SPLIT distance="625" swimtime="00:06:52.55" />
                    <SPLIT distance="650" swimtime="00:07:09.31" />
                    <SPLIT distance="675" swimtime="00:07:26.01" />
                    <SPLIT distance="700" swimtime="00:07:43.05" />
                    <SPLIT distance="725" swimtime="00:07:59.34" />
                    <SPLIT distance="750" swimtime="00:08:16.00" />
                    <SPLIT distance="775" swimtime="00:08:32.40" />
                    <SPLIT distance="800" swimtime="00:08:49.22" />
                    <SPLIT distance="825" swimtime="00:09:05.70" />
                    <SPLIT distance="850" swimtime="00:09:22.50" />
                    <SPLIT distance="875" swimtime="00:09:39.21" />
                    <SPLIT distance="900" swimtime="00:09:56.04" />
                    <SPLIT distance="925" swimtime="00:10:12.67" />
                    <SPLIT distance="950" swimtime="00:10:29.49" />
                    <SPLIT distance="975" swimtime="00:10:45.95" />
                    <SPLIT distance="1000" swimtime="00:11:02.71" />
                    <SPLIT distance="1025" swimtime="00:11:19.35" />
                    <SPLIT distance="1050" swimtime="00:11:36.12" />
                    <SPLIT distance="1075" swimtime="00:11:52.86" />
                    <SPLIT distance="1100" swimtime="00:12:09.47" />
                    <SPLIT distance="1125" swimtime="00:12:26.14" />
                    <SPLIT distance="1150" swimtime="00:12:43.05" />
                    <SPLIT distance="1175" swimtime="00:12:59.73" />
                    <SPLIT distance="1200" swimtime="00:13:16.48" />
                    <SPLIT distance="1225" swimtime="00:13:33.21" />
                    <SPLIT distance="1250" swimtime="00:13:49.99" />
                    <SPLIT distance="1275" swimtime="00:14:06.73" />
                    <SPLIT distance="1300" swimtime="00:14:23.35" />
                    <SPLIT distance="1325" swimtime="00:14:40.12" />
                    <SPLIT distance="1350" swimtime="00:14:56.97" />
                    <SPLIT distance="1375" swimtime="00:15:13.68" />
                    <SPLIT distance="1400" swimtime="00:15:30.53" />
                    <SPLIT distance="1425" swimtime="00:15:46.87" />
                    <SPLIT distance="1450" swimtime="00:16:03.64" />
                    <SPLIT distance="1475" swimtime="00:16:19.98" />
                    <SPLIT distance="1500" swimtime="00:16:35.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="South Africa">
              <RESULTS>
                <RESULT eventid="9" place="13" lane="7" heat="2" swimtime="00:03:25.51" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.80" />
                    <SPLIT distance="50" swimtime="00:00:22.97" />
                    <SPLIT distance="75" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:00:48.75" />
                    <SPLIT distance="125" swimtime="00:00:59.62" />
                    <SPLIT distance="150" swimtime="00:01:12.20" />
                    <SPLIT distance="175" swimtime="00:01:25.03" />
                    <SPLIT distance="200" swimtime="00:01:37.50" />
                    <SPLIT distance="225" swimtime="00:01:48.95" />
                    <SPLIT distance="250" swimtime="00:02:01.59" />
                    <SPLIT distance="275" swimtime="00:02:14.80" />
                    <SPLIT distance="300" swimtime="00:02:28.20" />
                    <SPLIT distance="325" swimtime="00:02:41.15" />
                    <SPLIT distance="350" swimtime="00:02:55.79" />
                    <SPLIT distance="375" swimtime="00:03:10.82" />
                    <SPLIT distance="400" swimtime="00:03:25.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="212656" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="108867" reactiontime="+26" />
                    <RELAYPOSITION number="3" athleteid="197938" reactiontime="+53" />
                    <RELAYPOSITION number="4" athleteid="154863" reactiontime="+76" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="South Africa">
              <RESULTS>
                <RESULT eventid="26" place="12" lane="8" heat="1" swimtime="00:01:29.27" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.59" />
                    <SPLIT distance="50" swimtime="00:00:21.84" />
                    <SPLIT distance="75" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:00:44.09" />
                    <SPLIT distance="125" swimtime="00:00:55.33" />
                    <SPLIT distance="150" swimtime="00:01:07.52" />
                    <SPLIT distance="175" swimtime="00:01:18.12" />
                    <SPLIT distance="200" swimtime="00:01:29.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="108867" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="212656" reactiontime="+26" />
                    <RELAYPOSITION number="3" athleteid="197938" reactiontime="+47" />
                    <RELAYPOSITION number="4" athleteid="170357" reactiontime="+59" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="South Africa">
              <RESULTS>
                <RESULT eventid="27" place="11" lane="3" heat="2" swimtime="00:01:33.28" reactiontime="+66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:21.83" />
                    <SPLIT distance="75" swimtime="00:00:32.06" />
                    <SPLIT distance="100" swimtime="00:00:43.67" />
                    <SPLIT distance="125" swimtime="00:00:55.07" />
                    <SPLIT distance="150" swimtime="00:01:07.96" />
                    <SPLIT distance="175" swimtime="00:01:20.18" />
                    <SPLIT distance="200" swimtime="00:01:33.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="108867" reactiontime="+66" />
                    <RELAYPOSITION number="2" athleteid="212656" reactiontime="+7" />
                    <RELAYPOSITION number="3" athleteid="191644" reactiontime="+11" />
                    <RELAYPOSITION number="4" athleteid="210937" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="South Africa">
              <RESULTS>
                <RESULT eventid="8" place="13" lane="2" heat="1" swimtime="00:03:41.57" reactiontime="+78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.05" />
                    <SPLIT distance="50" swimtime="00:00:27.20" />
                    <SPLIT distance="75" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:00:56.97" />
                    <SPLIT distance="125" swimtime="00:01:08.45" />
                    <SPLIT distance="150" swimtime="00:01:21.91" />
                    <SPLIT distance="175" swimtime="00:01:36.02" />
                    <SPLIT distance="200" swimtime="00:01:50.30" />
                    <SPLIT distance="225" swimtime="00:02:03.10" />
                    <SPLIT distance="250" swimtime="00:02:17.47" />
                    <SPLIT distance="275" swimtime="00:02:32.39" />
                    <SPLIT distance="300" swimtime="00:02:47.38" />
                    <SPLIT distance="325" swimtime="00:02:59.51" />
                    <SPLIT distance="350" swimtime="00:03:13.43" />
                    <SPLIT distance="375" swimtime="00:03:27.59" />
                    <SPLIT distance="400" swimtime="00:03:41.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="210937" reactiontime="+78" />
                    <RELAYPOSITION number="2" athleteid="191644" reactiontime="-2" />
                    <RELAYPOSITION number="3" athleteid="108899" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="144092" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="South Africa">
              <RESULTS>
                <RESULT eventid="47" place="12" lane="7" heat="2" swimtime="00:03:59.64" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.43" />
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="75" swimtime="00:00:45.09" />
                    <SPLIT distance="100" swimtime="00:01:00.30" />
                    <SPLIT distance="125" swimtime="00:01:14.95" />
                    <SPLIT distance="150" swimtime="00:01:32.08" />
                    <SPLIT distance="175" swimtime="00:01:49.61" />
                    <SPLIT distance="200" swimtime="00:02:07.70" />
                    <SPLIT distance="225" swimtime="00:02:19.59" />
                    <SPLIT distance="250" swimtime="00:02:34.19" />
                    <SPLIT distance="275" swimtime="00:02:49.62" />
                    <SPLIT distance="300" swimtime="00:03:05.38" />
                    <SPLIT distance="325" swimtime="00:03:17.12" />
                    <SPLIT distance="350" swimtime="00:03:30.95" />
                    <SPLIT distance="375" swimtime="00:03:45.15" />
                    <SPLIT distance="400" swimtime="00:03:59.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="210937" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="108899" reactiontime="+45" />
                    <RELAYPOSITION number="3" athleteid="144092" reactiontime="+44" />
                    <RELAYPOSITION number="4" athleteid="191644" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="South Africa">
              <RESULTS>
                <RESULT eventid="17" place="10" lane="2" heat="1" swimtime="00:08:04.85" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="75" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:01.29" />
                    <SPLIT distance="125" swimtime="00:01:16.56" />
                    <SPLIT distance="150" swimtime="00:01:32.20" />
                    <SPLIT distance="175" swimtime="00:01:47.64" />
                    <SPLIT distance="200" swimtime="00:02:02.67" />
                    <SPLIT distance="225" swimtime="00:02:15.68" />
                    <SPLIT distance="250" swimtime="00:02:30.44" />
                    <SPLIT distance="275" swimtime="00:02:45.51" />
                    <SPLIT distance="300" swimtime="00:03:00.82" />
                    <SPLIT distance="325" swimtime="00:03:16.44" />
                    <SPLIT distance="350" swimtime="00:03:32.44" />
                    <SPLIT distance="375" swimtime="00:03:48.64" />
                    <SPLIT distance="400" swimtime="00:04:04.44" />
                    <SPLIT distance="425" swimtime="00:04:17.72" />
                    <SPLIT distance="450" swimtime="00:04:32.52" />
                    <SPLIT distance="475" swimtime="00:04:47.60" />
                    <SPLIT distance="500" swimtime="00:05:03.05" />
                    <SPLIT distance="525" swimtime="00:05:18.98" />
                    <SPLIT distance="550" swimtime="00:05:35.19" />
                    <SPLIT distance="575" swimtime="00:05:51.40" />
                    <SPLIT distance="600" swimtime="00:06:07.18" />
                    <SPLIT distance="625" swimtime="00:06:19.36" />
                    <SPLIT distance="650" swimtime="00:06:33.62" />
                    <SPLIT distance="675" swimtime="00:06:48.38" />
                    <SPLIT distance="700" swimtime="00:07:03.40" />
                    <SPLIT distance="725" swimtime="00:07:18.61" />
                    <SPLIT distance="750" swimtime="00:07:34.15" />
                    <SPLIT distance="775" swimtime="00:07:49.69" />
                    <SPLIT distance="800" swimtime="00:08:04.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="170443" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="197620" reactiontime="+63" />
                    <RELAYPOSITION number="3" athleteid="108899" reactiontime="+44" />
                    <RELAYPOSITION number="4" athleteid="144092" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="South Africa">
              <RESULTS>
                <RESULT eventid="25" place="11" lane="2" heat="1" swimtime="00:01:40.80" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:24.33" />
                    <SPLIT distance="75" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:00:49.47" />
                    <SPLIT distance="125" swimtime="00:01:02.18" />
                    <SPLIT distance="150" swimtime="00:01:15.55" />
                    <SPLIT distance="175" swimtime="00:01:27.70" />
                    <SPLIT distance="200" swimtime="00:01:40.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="191644" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="144092" reactiontime="+42" />
                    <RELAYPOSITION number="3" athleteid="108899" reactiontime="+44" />
                    <RELAYPOSITION number="4" athleteid="210937" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="South Africa">
              <RESULTS>
                <RESULT eventid="34" place="13" lane="7" heat="2" swimtime="00:01:53.76" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                    <SPLIT distance="50" swimtime="00:00:28.24" />
                    <SPLIT distance="75" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:00:59.70" />
                    <SPLIT distance="125" swimtime="00:01:11.63" />
                    <SPLIT distance="150" swimtime="00:01:26.57" />
                    <SPLIT distance="175" swimtime="00:01:39.86" />
                    <SPLIT distance="200" swimtime="00:01:53.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="210937" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="108899" reactiontime="+46" />
                    <RELAYPOSITION number="3" athleteid="191644" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="170443" reactiontime="+68" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="South Africa">
              <RESULTS>
                <RESULT eventid="11" place="17" lane="3" heat="3" swimtime="00:01:43.07" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                    <SPLIT distance="75" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:00:55.73" />
                    <SPLIT distance="125" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:18.78" />
                    <SPLIT distance="175" swimtime="00:01:30.27" />
                    <SPLIT distance="200" swimtime="00:01:43.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="210937" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="212656" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="108867" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="191644" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="South Africa">
              <RESULTS>
                <RESULT eventid="35" place="14" lane="2" heat="2" swimtime="00:01:37.14" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:22.96" />
                    <SPLIT distance="75" swimtime="00:00:36.25" />
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                    <SPLIT distance="125" swimtime="00:01:02.16" />
                    <SPLIT distance="150" swimtime="00:01:14.86" />
                    <SPLIT distance="175" swimtime="00:01:25.53" />
                    <SPLIT distance="200" swimtime="00:01:37.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="170357" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="197938" reactiontime="+44" />
                    <RELAYPOSITION number="3" athleteid="108867" reactiontime="+47" />
                    <RELAYPOSITION number="4" athleteid="212656" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Russian Swimming Federation" shortname="RSF" code="RSF" nation="RSF" type="NOC">
          <ATHLETES />
        </CLUB>
        <CLUB name="Russian Federation" shortname="RUS" code="RUS" nation="RUS" type="NOC">
          <ATHLETES />
        </CLUB>
        <CLUB name="Rwanda" shortname="RWA" code="RWA" nation="RWA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="165326" lastname="NIYIBIZI" firstname="Cedrick" gender="M" birthdate="2001-01-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.44" eventid="14" heat="2" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.75" eventid="31" heat="3" lane="5">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="78" lane="3" heat="2" heatid="20014" swimtime="00:00:55.87" reactiontime="+71" points="516">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.37" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                    <SPLIT distance="75" swimtime="00:00:41.09" />
                    <SPLIT distance="100" swimtime="00:00:55.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="64" lane="5" heat="3" heatid="30031" swimtime="00:00:24.95" reactiontime="+69" points="527">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:24.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Samoa" shortname="SAM" code="SAM" nation="SAM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="100651" lastname="SCHUSTER" firstname="Brandon" gender="M" birthdate="1998-04-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.72" eventid="16" heat="2" lane="1">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.56" eventid="31" heat="3" lane="4">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="51" lane="1" heat="2" heatid="20016" swimtime="00:01:01.96" reactiontime="+64" points="710">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.29" />
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                    <SPLIT distance="75" swimtime="00:00:45.13" />
                    <SPLIT distance="100" swimtime="00:01:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="55" lane="4" heat="3" heatid="30031" swimtime="00:00:23.71" reactiontime="+66" points="614">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196120" lastname="FROST" firstname="Kokoro" gender="M" birthdate="2002-09-14">
              <ENTRIES>
                <ENTRY entrytime="00:00:26.44" eventid="19" heat="1" lane="5">
                  <MEETINFO date="2022-08-26" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.08" eventid="5" heat="4" lane="8">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="37" lane="5" heat="1" heatid="10019" swimtime="00:00:26.18" reactiontime="+59" points="611">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.66" />
                    <SPLIT distance="50" swimtime="00:00:26.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="53" lane="8" heat="4" heatid="40005" swimtime="00:00:25.03" reactiontime="+63" points="656">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:25.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201156" lastname="BORG" firstname="Olivia" gender="F" birthdate="2001-01-19">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:01.13" eventid="38" heat="1" lane="5">
                  <MEETINFO date="2022-05-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.37" eventid="4" heat="3" lane="3">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="25" lane="5" heat="1" heatid="10038" swimtime="00:01:00.13" reactiontime="+71" points="748">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                    <SPLIT distance="75" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:01:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="28" lane="3" heat="3" heatid="30004" swimtime="00:00:27.09" reactiontime="+75" points="728">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.57" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213131" lastname="BROWN" firstname="Kaiya" gender="F" birthdate="2004-04-17">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:01.83" eventid="13" heat="3" lane="3">
                  <MEETINFO date="2022-08-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.84" eventid="30" heat="3" lane="5">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="49" lane="3" heat="3" heatid="30013" swimtime="00:00:59.17" reactiontime="+69" points="612">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="75" swimtime="00:00:43.71" />
                    <SPLIT distance="100" swimtime="00:00:59.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="40" lane="5" heat="3" heatid="30030" swimtime="00:00:27.43" reactiontime="+70" points="584">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Samoa">
              <RESULTS>
                <RESULT eventid="27" place="19" lane="8" heat="3" swimtime="00:01:39.49" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:24.02" />
                    <SPLIT distance="75" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:00:47.04" />
                    <SPLIT distance="125" swimtime="00:00:59.99" />
                    <SPLIT distance="150" swimtime="00:01:14.10" />
                    <SPLIT distance="175" swimtime="00:01:26.10" />
                    <SPLIT distance="200" swimtime="00:01:39.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196120" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="100651" reactiontime="+26" />
                    <RELAYPOSITION number="3" athleteid="213131" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="201156" reactiontime="+28" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Samoa">
              <RESULTS>
                <RESULT eventid="11" place="23" lane="8" heat="3" swimtime="00:01:47.91" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                    <SPLIT distance="75" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:00:54.08" />
                    <SPLIT distance="125" swimtime="00:01:06.41" />
                    <SPLIT distance="150" swimtime="00:01:21.14" />
                    <SPLIT distance="175" swimtime="00:01:33.99" />
                    <SPLIT distance="200" swimtime="00:01:47.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="196120" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="100651" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="201156" reactiontime="+47" />
                    <RELAYPOSITION number="4" athleteid="213131" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Senegal" shortname="SEN" code="SEN" nation="SEN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="166107" lastname="AIMABLE" firstname="Steven" gender="M" birthdate="1999-02-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.64" eventid="39" heat="3" lane="4">
                  <MEETINFO date="2021-07-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.08" eventid="31" heat="5" lane="6">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="37" lane="4" heat="3" heatid="30039" swimtime="00:00:53.08" reactiontime="+58" points="729">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.24" />
                    <SPLIT distance="50" swimtime="00:00:24.73" />
                    <SPLIT distance="75" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:00:53.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="48" lane="6" heat="5" heatid="50031" swimtime="00:00:22.42" reactiontime="+59" points="727">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.85" />
                    <SPLIT distance="50" swimtime="00:00:22.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198110" lastname="DIOP" firstname="Oumy" gender="F" birthdate="2003-08-29">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.24" eventid="38" heat="1" lane="3">
                  <MEETINFO date="2022-08-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:58.33" eventid="13" heat="4" lane="3">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="27" lane="3" heat="1" heatid="10038" swimtime="00:01:01.54" reactiontime="+71" points="698">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:28.69" />
                    <SPLIT distance="75" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="46" lane="3" heat="4" heatid="40013" swimtime="00:00:58.47" reactiontime="+70" points="634">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                    <SPLIT distance="75" swimtime="00:00:43.04" />
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Singapore" shortname="SGP" code="SGP" nation="SGP" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="129524" lastname="ANG" firstname="Maximillian Wei" gender="M" birthdate="2001-03-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.72" eventid="16" heat="5" lane="1">
                  <MEETINFO date="2021-11-26" />
                </ENTRY>
                <ENTRY entrytime="00:02:08.49" eventid="29" heat="3" lane="8">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="00:01:57.18" eventid="7" heat="3" lane="1">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.23" eventid="41" heat="4" lane="6">
                  <MEETINFO date="2022-08-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.47" eventid="23" heat="2" lane="5">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="22" lane="1" heat="5" heatid="50016" swimtime="00:00:58.10" reactiontime="+63" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                    <SPLIT distance="75" swimtime="00:00:42.51" />
                    <SPLIT distance="100" swimtime="00:00:58.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="19" lane="8" heat="3" heatid="30029" swimtime="00:02:08.12" reactiontime="+72" points="824">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="75" swimtime="00:00:45.04" />
                    <SPLIT distance="100" swimtime="00:01:01.45" />
                    <SPLIT distance="125" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:01:34.65" />
                    <SPLIT distance="175" swimtime="00:01:51.26" />
                    <SPLIT distance="200" swimtime="00:02:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="28" lane="1" heat="3" heatid="30007" swimtime="00:01:59.11" reactiontime="+64" points="779">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.32" />
                    <SPLIT distance="50" swimtime="00:00:25.21" />
                    <SPLIT distance="75" swimtime="00:00:40.93" />
                    <SPLIT distance="100" swimtime="00:00:55.78" />
                    <SPLIT distance="125" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:29.56" />
                    <SPLIT distance="175" swimtime="00:01:45.14" />
                    <SPLIT distance="200" swimtime="00:01:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="28" lane="6" heat="4" heatid="40041" swimtime="00:00:27.09" reactiontime="+62" points="781">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="29" lane="5" heat="2" heatid="20023" swimtime="00:00:54.79" reactiontime="+62" points="727">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.27" />
                    <SPLIT distance="50" swimtime="00:00:25.34" />
                    <SPLIT distance="75" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:00:54.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124017" lastname="TEONG" firstname="Tzen Wei" gender="M" birthdate="1997-10-17">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.88" eventid="39">
                  <MEETINFO date="2021-11-26" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.24" eventid="5" heat="10" lane="3">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.27" eventid="31" heat="10" lane="7">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="105" place="4" lane="1" heat="1" heatid="10105" swimtime="00:00:22.01" reactiontime="+58" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.92" />
                    <SPLIT distance="50" swimtime="00:00:22.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="1" lane="3" heat="10" heatid="100005" swimtime="00:00:22.01" reactiontime="+62" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.98" />
                    <SPLIT distance="50" swimtime="00:00:22.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="7" lane="4" heat="1" heatid="10205" swimtime="00:00:22.18" reactiontime="+59" points="942">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.07" />
                    <SPLIT distance="50" swimtime="00:00:22.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="17" lane="7" heat="10" heatid="100031" swimtime="00:00:21.30" reactiontime="+61" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.12" />
                    <SPLIT distance="50" swimtime="00:00:21.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="11" lane="8" heat="1" heatid="10231" swimtime="00:00:21.09" reactiontime="+60" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.12" />
                    <SPLIT distance="50" swimtime="00:00:21.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197628" lastname="SIM" firstname="En Yi Letitia" gender="F" birthdate="2003-03-03">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.44" eventid="15" heat="6" lane="1">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:27.44" eventid="28" heat="2" lane="7">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.30" eventid="6" heat="2" lane="8">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.75" eventid="40" heat="4" lane="4">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="28" lane="1" heat="6" heatid="60015" swimtime="00:01:06.49" reactiontime="+65" points="824">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.32" />
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="75" swimtime="00:00:48.65" />
                    <SPLIT distance="100" swimtime="00:01:06.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="14" lane="7" heat="2" heatid="20028" swimtime="00:02:21.60" reactiontime="+65" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="75" swimtime="00:00:50.21" />
                    <SPLIT distance="100" swimtime="00:01:08.28" />
                    <SPLIT distance="125" swimtime="00:01:26.21" />
                    <SPLIT distance="150" swimtime="00:01:44.29" />
                    <SPLIT distance="175" swimtime="00:02:02.89" />
                    <SPLIT distance="200" swimtime="00:02:21.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="18" lane="8" heat="2" heatid="20006" swimtime="00:02:09.82" reactiontime="+65" points="827">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.69" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="75" swimtime="00:00:45.13" />
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                    <SPLIT distance="125" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:01:38.39" />
                    <SPLIT distance="175" swimtime="00:01:54.70" />
                    <SPLIT distance="200" swimtime="00:02:09.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="22" lane="4" heat="4" heatid="40040" swimtime="00:00:30.59" reactiontime="+62" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129528" lastname="GAN" firstname="Ching Hwee" gender="F" birthdate="2003-07-22">
              <ENTRIES>
                <ENTRY entrytime="00:01:58.85" eventid="43" heat="4" lane="8">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:04:07.50" eventid="1" heat="2" lane="5">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:08:22.91" eventid="12" heat="0" lane="-1">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:16:32.43" eventid="33" heat="2" lane="2">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="-1" lane="8" heat="4" heatid="40043" swimtime="NT" status="DNS" />
                <RESULT eventid="1" place="-1" lane="5" heat="2" heatid="20001" swimtime="NT" status="DNS" />
                <RESULT eventid="112" place="-1" lane="1" heat="5" heatid="30112" swimtime="NT" status="DNS" />
                <RESULT eventid="133" place="-1" lane="2" heat="2" heatid="20033" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Saint Kitts &amp; Nevis" shortname="SKN" code="SKN" nation="SKN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="163124" lastname="HARDING-MARLIN" firstname="Jennifer Lynn" gender="F" birthdate="1992-06-11">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="45" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="22" heat="1" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="34" lane="3" heat="1" heatid="10045" swimtime="00:02:31.55" reactiontime="+75" points="483">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="75" swimtime="00:00:53.09" />
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                    <SPLIT distance="125" swimtime="00:01:32.22" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                    <SPLIT distance="175" swimtime="00:02:12.47" />
                    <SPLIT distance="200" swimtime="00:02:31.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="28" lane="2" heat="1" heatid="10022" swimtime="00:01:13.46" reactiontime="+78" points="455">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.13" />
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="75" swimtime="00:00:55.59" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Sierra Leone" shortname="SLE" code="SLE" nation="SLE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="201909" lastname="KAMARA" firstname="Sheku" gender="M" birthdate="1999-11-19">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="19" heat="1" lane="2" />
                <ENTRY entrytime="NT" eventid="41" heat="2" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="-1" lane="2" heat="1" heatid="10019" swimtime="NT" status="DNS" />
                <RESULT eventid="41" place="-1" lane="2" heat="2" heatid="20041" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150000" lastname="BANGURA" firstname="Sheku" gender="M" birthdate="2003-04-15">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5" heat="2" lane="7" />
                <ENTRY entrytime="00:00:29.90" eventid="31" heat="2" lane="6">
                  <MEETINFO date="2021-10-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="-1" lane="7" heat="2" heatid="20005" swimtime="NT" status="DNS" />
                <RESULT eventid="31" place="77" lane="6" heat="2" heatid="20031" swimtime="00:00:29.38" reactiontime="+68" points="323">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198079" lastname="YONGAI" firstname="Mary" gender="F" birthdate="2003-03-13">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="40" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="43" lane="4" heat="1" heatid="10040" swimtime="00:00:46.98" reactiontime="+75" points="224">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.99" />
                    <SPLIT distance="50" swimtime="00:00:46.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="58" lane="1" heat="1" heatid="10030" swimtime="00:00:41.41" reactiontime="+84" points="169">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.65" />
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214442" lastname="KAMARA" firstname="Yaba" gender="F" birthdate="2006-01-27">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="4" heat="1" lane="5" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="-1" lane="5" heat="1" heatid="10004" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Slovenia" shortname="SLO" code="SLO" nation="SLO" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="108709" lastname="STEVENS" firstname="Peter " gender="M" birthdate="1995-06-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.92" eventid="16" heat="6" lane="8">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.10" eventid="41" heat="9" lane="3">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="27" lane="8" heat="6" heatid="60016" swimtime="00:00:58.31" reactiontime="+62" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.10" />
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                    <SPLIT distance="75" swimtime="00:00:42.38" />
                    <SPLIT distance="100" swimtime="00:00:58.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="10" lane="3" heat="9" heatid="90041" swimtime="00:00:26.31" reactiontime="+59" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.87" />
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="13" lane="2" heat="1" heatid="10241" swimtime="00:00:26.33" reactiontime="+60" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:26.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122192" lastname="VOVK" firstname="Tara" gender="F" birthdate="2000-02-15">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="15" heat="1" lane="1" />
                <ENTRY entrytime="00:00:31.12" eventid="40" heat="4" lane="2">
                  <MEETINFO date="2022-03-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="26" lane="1" heat="1" heatid="10015" swimtime="00:01:06.29" reactiontime="+71" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="75" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="19" lane="2" heat="4" heatid="40040" swimtime="00:00:30.39" reactiontime="+60" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122197" lastname="KLANCAR" firstname="Neza" gender="F" birthdate="2000-02-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:54.24" eventid="13" heat="6" lane="5">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.50" eventid="4" heat="6" lane="8">
                  <MEETINFO date="2022-07-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.96" eventid="30" heat="8" lane="8">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:00.87" eventid="22" heat="3" lane="1">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="22" lane="5" heat="6" heatid="60013" swimtime="00:00:53.81" reactiontime="+66" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.38" />
                    <SPLIT distance="50" swimtime="00:00:25.87" />
                    <SPLIT distance="75" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:00:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="17" lane="8" heat="6" heatid="60004" swimtime="00:00:25.85" reactiontime="+66" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="304" place="18" lane="4" heat="1" heatid="10304" swimtime="00:00:25.85" reactiontime="+65" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="9" lane="8" heat="8" heatid="80030" swimtime="00:00:24.16" reactiontime="+67" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:24.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="9" lane="2" heat="2" heatid="20230" swimtime="00:00:24.13" reactiontime="+67" points="858">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="9" lane="1" heat="3" heatid="30022" swimtime="00:00:59.42" reactiontime="+68" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:27.21" />
                    <SPLIT distance="75" swimtime="00:00:44.96" />
                    <SPLIT distance="100" swimtime="00:00:59.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="9" lane="2" heat="2" heatid="20222" swimtime="00:00:59.27" reactiontime="+71" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:27.17" />
                    <SPLIT distance="75" swimtime="00:00:44.67" />
                    <SPLIT distance="100" swimtime="00:00:59.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="140817" lastname="FAIN" firstname="Katja" gender="F" birthdate="2001-08-31">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.48" eventid="43" heat="3" lane="3">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:04:03.52" eventid="1" heat="3" lane="7">
                  <MEETINFO date="2021-10-07" />
                </ENTRY>
                <ENTRY entrytime="00:16:13.42" eventid="33" heat="2" lane="4">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="10" lane="3" heat="3" heatid="30043" swimtime="00:01:54.96" reactiontime="+73" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:42.06" />
                    <SPLIT distance="100" swimtime="00:00:56.77" />
                    <SPLIT distance="125" swimtime="00:01:11.31" />
                    <SPLIT distance="150" swimtime="00:01:26.02" />
                    <SPLIT distance="175" swimtime="00:01:40.82" />
                    <SPLIT distance="200" swimtime="00:01:54.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="101" place="5" lane="1" heat="1" heatid="10101" swimtime="00:04:01.46" reactiontime="+71" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="75" swimtime="00:00:43.24" />
                    <SPLIT distance="100" swimtime="00:00:58.59" />
                    <SPLIT distance="125" swimtime="00:01:13.89" />
                    <SPLIT distance="150" swimtime="00:01:29.20" />
                    <SPLIT distance="175" swimtime="00:01:44.64" />
                    <SPLIT distance="200" swimtime="00:02:00.07" />
                    <SPLIT distance="225" swimtime="00:02:15.49" />
                    <SPLIT distance="250" swimtime="00:02:31.01" />
                    <SPLIT distance="275" swimtime="00:02:46.42" />
                    <SPLIT distance="300" swimtime="00:03:01.78" />
                    <SPLIT distance="325" swimtime="00:03:17.20" />
                    <SPLIT distance="350" swimtime="00:03:32.43" />
                    <SPLIT distance="375" swimtime="00:03:47.49" />
                    <SPLIT distance="400" swimtime="00:04:01.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="7" lane="7" heat="3" heatid="30001" swimtime="00:04:02.13" reactiontime="+73" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="75" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:00:58.77" />
                    <SPLIT distance="125" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:29.51" />
                    <SPLIT distance="175" swimtime="00:01:44.65" />
                    <SPLIT distance="200" swimtime="00:02:00.26" />
                    <SPLIT distance="225" swimtime="00:02:15.62" />
                    <SPLIT distance="250" swimtime="00:02:30.92" />
                    <SPLIT distance="275" swimtime="00:02:46.42" />
                    <SPLIT distance="300" swimtime="00:03:01.97" />
                    <SPLIT distance="325" swimtime="00:03:17.10" />
                    <SPLIT distance="350" swimtime="00:03:32.54" />
                    <SPLIT distance="375" swimtime="00:03:47.84" />
                    <SPLIT distance="400" swimtime="00:04:02.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="9" lane="4" heat="2" heatid="20033" swimtime="00:16:12.06" reactiontime="+72" points="842">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="75" swimtime="00:00:45.06" />
                    <SPLIT distance="100" swimtime="00:01:00.68" />
                    <SPLIT distance="125" swimtime="00:01:16.62" />
                    <SPLIT distance="150" swimtime="00:01:32.51" />
                    <SPLIT distance="175" swimtime="00:01:48.39" />
                    <SPLIT distance="200" swimtime="00:02:04.31" />
                    <SPLIT distance="225" swimtime="00:02:20.22" />
                    <SPLIT distance="250" swimtime="00:02:36.44" />
                    <SPLIT distance="275" swimtime="00:02:52.59" />
                    <SPLIT distance="300" swimtime="00:03:08.69" />
                    <SPLIT distance="325" swimtime="00:03:24.74" />
                    <SPLIT distance="350" swimtime="00:03:40.74" />
                    <SPLIT distance="375" swimtime="00:03:56.89" />
                    <SPLIT distance="400" swimtime="00:04:13.04" />
                    <SPLIT distance="425" swimtime="00:04:29.15" />
                    <SPLIT distance="450" swimtime="00:04:45.30" />
                    <SPLIT distance="475" swimtime="00:05:01.46" />
                    <SPLIT distance="500" swimtime="00:05:17.54" />
                    <SPLIT distance="525" swimtime="00:05:33.56" />
                    <SPLIT distance="550" swimtime="00:05:49.63" />
                    <SPLIT distance="575" swimtime="00:06:05.90" />
                    <SPLIT distance="600" swimtime="00:06:22.06" />
                    <SPLIT distance="625" swimtime="00:06:38.33" />
                    <SPLIT distance="650" swimtime="00:06:54.57" />
                    <SPLIT distance="675" swimtime="00:07:10.87" />
                    <SPLIT distance="700" swimtime="00:07:27.06" />
                    <SPLIT distance="725" swimtime="00:07:43.28" />
                    <SPLIT distance="750" swimtime="00:07:59.58" />
                    <SPLIT distance="775" swimtime="00:08:15.82" />
                    <SPLIT distance="800" swimtime="00:08:32.09" />
                    <SPLIT distance="825" swimtime="00:08:48.42" />
                    <SPLIT distance="850" swimtime="00:09:04.87" />
                    <SPLIT distance="875" swimtime="00:09:21.10" />
                    <SPLIT distance="900" swimtime="00:09:37.42" />
                    <SPLIT distance="925" swimtime="00:09:53.84" />
                    <SPLIT distance="950" swimtime="00:10:10.18" />
                    <SPLIT distance="975" swimtime="00:10:26.74" />
                    <SPLIT distance="1000" swimtime="00:10:43.41" />
                    <SPLIT distance="1025" swimtime="00:10:59.91" />
                    <SPLIT distance="1050" swimtime="00:11:16.54" />
                    <SPLIT distance="1075" swimtime="00:11:33.17" />
                    <SPLIT distance="1100" swimtime="00:11:49.78" />
                    <SPLIT distance="1125" swimtime="00:12:06.43" />
                    <SPLIT distance="1150" swimtime="00:12:23.09" />
                    <SPLIT distance="1175" swimtime="00:12:39.88" />
                    <SPLIT distance="1200" swimtime="00:12:56.54" />
                    <SPLIT distance="1225" swimtime="00:13:13.07" />
                    <SPLIT distance="1250" swimtime="00:13:29.72" />
                    <SPLIT distance="1275" swimtime="00:13:46.25" />
                    <SPLIT distance="1300" swimtime="00:14:02.71" />
                    <SPLIT distance="1325" swimtime="00:14:19.23" />
                    <SPLIT distance="1350" swimtime="00:14:35.85" />
                    <SPLIT distance="1375" swimtime="00:14:52.15" />
                    <SPLIT distance="1400" swimtime="00:15:08.48" />
                    <SPLIT distance="1425" swimtime="00:15:24.79" />
                    <SPLIT distance="1450" swimtime="00:15:40.98" />
                    <SPLIT distance="1475" swimtime="00:15:57.00" />
                    <SPLIT distance="1500" swimtime="00:16:12.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Suspended Member Federation" shortname="SMF" code="SMF" nation="SMF" type="">
          <ATHLETES>
            <ATHLETE athleteid="201883" lastname="HART" firstname="Ivan" gender="M" birthdate="2006-09-22">
              <ENTRIES>
                <ENTRY entrytime="00:16:45.33" eventid="10" heat="1" lane="3">
                  <MEETINFO date="2022-04-07" />
                </ENTRY>
                <ENTRY entrytime="00:04:15.40" eventid="24" heat="1" lane="2">
                  <MEETINFO date="2022-04-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="16" lane="3" heat="1" heatid="10010" swimtime="00:16:07.94" reactiontime="+72" points="669">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="75" swimtime="00:00:44.11" />
                    <SPLIT distance="100" swimtime="00:00:59.71" />
                    <SPLIT distance="125" swimtime="00:01:15.69" />
                    <SPLIT distance="150" swimtime="00:01:31.61" />
                    <SPLIT distance="175" swimtime="00:01:47.55" />
                    <SPLIT distance="200" swimtime="00:02:03.30" />
                    <SPLIT distance="225" swimtime="00:02:19.16" />
                    <SPLIT distance="250" swimtime="00:02:35.14" />
                    <SPLIT distance="275" swimtime="00:02:51.09" />
                    <SPLIT distance="300" swimtime="00:03:07.04" />
                    <SPLIT distance="325" swimtime="00:03:22.90" />
                    <SPLIT distance="350" swimtime="00:03:38.88" />
                    <SPLIT distance="375" swimtime="00:03:54.92" />
                    <SPLIT distance="400" swimtime="00:04:11.11" />
                    <SPLIT distance="425" swimtime="00:04:27.18" />
                    <SPLIT distance="450" swimtime="00:04:43.24" />
                    <SPLIT distance="475" swimtime="00:04:59.36" />
                    <SPLIT distance="500" swimtime="00:05:15.63" />
                    <SPLIT distance="525" swimtime="00:05:31.87" />
                    <SPLIT distance="550" swimtime="00:05:48.03" />
                    <SPLIT distance="575" swimtime="00:06:04.28" />
                    <SPLIT distance="600" swimtime="00:06:20.77" />
                    <SPLIT distance="625" swimtime="00:06:36.94" />
                    <SPLIT distance="650" swimtime="00:06:53.35" />
                    <SPLIT distance="675" swimtime="00:07:09.27" />
                    <SPLIT distance="700" swimtime="00:07:25.57" />
                    <SPLIT distance="725" swimtime="00:07:41.78" />
                    <SPLIT distance="750" swimtime="00:07:58.11" />
                    <SPLIT distance="775" swimtime="00:08:14.26" />
                    <SPLIT distance="800" swimtime="00:08:30.53" />
                    <SPLIT distance="825" swimtime="00:08:46.72" />
                    <SPLIT distance="850" swimtime="00:09:02.91" />
                    <SPLIT distance="875" swimtime="00:09:19.21" />
                    <SPLIT distance="900" swimtime="00:09:35.71" />
                    <SPLIT distance="925" swimtime="00:09:52.11" />
                    <SPLIT distance="950" swimtime="00:10:08.50" />
                    <SPLIT distance="975" swimtime="00:10:25.04" />
                    <SPLIT distance="1000" swimtime="00:10:41.53" />
                    <SPLIT distance="1025" swimtime="00:10:58.03" />
                    <SPLIT distance="1050" swimtime="00:11:14.47" />
                    <SPLIT distance="1075" swimtime="00:11:30.72" />
                    <SPLIT distance="1100" swimtime="00:11:47.17" />
                    <SPLIT distance="1125" swimtime="00:12:03.56" />
                    <SPLIT distance="1150" swimtime="00:12:20.02" />
                    <SPLIT distance="1175" swimtime="00:12:36.48" />
                    <SPLIT distance="1200" swimtime="00:12:52.96" />
                    <SPLIT distance="1225" swimtime="00:13:09.30" />
                    <SPLIT distance="1250" swimtime="00:13:25.53" />
                    <SPLIT distance="1275" swimtime="00:13:41.81" />
                    <SPLIT distance="1300" swimtime="00:13:58.31" />
                    <SPLIT distance="1325" swimtime="00:14:14.81" />
                    <SPLIT distance="1350" swimtime="00:14:31.18" />
                    <SPLIT distance="1375" swimtime="00:14:47.40" />
                    <SPLIT distance="1400" swimtime="00:15:03.96" />
                    <SPLIT distance="1425" swimtime="00:15:20.16" />
                    <SPLIT distance="1450" swimtime="00:15:36.45" />
                    <SPLIT distance="1475" swimtime="00:15:52.55" />
                    <SPLIT distance="1500" swimtime="00:16:07.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="33" lane="2" heat="1" heatid="10024" swimtime="00:04:08.64" reactiontime="+63" points="622">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:00:57.67" />
                    <SPLIT distance="125" swimtime="00:01:13.12" />
                    <SPLIT distance="150" swimtime="00:01:28.83" />
                    <SPLIT distance="175" swimtime="00:01:44.60" />
                    <SPLIT distance="200" swimtime="00:02:00.69" />
                    <SPLIT distance="225" swimtime="00:02:16.67" />
                    <SPLIT distance="250" swimtime="00:02:32.76" />
                    <SPLIT distance="275" swimtime="00:02:48.70" />
                    <SPLIT distance="300" swimtime="00:03:05.13" />
                    <SPLIT distance="325" swimtime="00:03:21.53" />
                    <SPLIT distance="350" swimtime="00:03:37.81" />
                    <SPLIT distance="375" swimtime="00:03:53.76" />
                    <SPLIT distance="400" swimtime="00:04:08.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214452" lastname="MURAVVEJ" firstname="Aryen" gender="M" birthdate="2005-05-11">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="5" heat="1" lane="4" />
                <ENTRY entrytime="NT" eventid="31" heat="1" lane="3" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="56" lane="4" heat="1" heatid="10005" swimtime="00:00:26.59" reactiontime="+59" points="547">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.44" />
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="56" lane="3" heat="1" heatid="10031" swimtime="00:00:24.08" reactiontime="+57" points="586">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:24.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130798" lastname="THORPE" firstname="Imara Bella Patricia" gender="F" birthdate="2001-02-20">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.16" eventid="38" heat="1" lane="2">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.78" eventid="4" heat="3" lane="2">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="28" lane="2" heat="1" heatid="10038" swimtime="00:01:01.84" reactiontime="+61" points="687">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                    <SPLIT distance="75" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:01.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="29" lane="2" heat="3" heatid="30004" swimtime="00:00:27.38" reactiontime="+60" points="705">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:27.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201886" lastname="ALI" firstname="Lubaina" gender="F" birthdate="2005-12-18">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.74" eventid="13" heat="3" lane="7">
                  <MEETINFO date="2021-10-11" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.19" eventid="43" heat="1" lane="6">
                  <MEETINFO date="2021-10-12" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="53" lane="7" heat="3" heatid="30013" swimtime="00:01:00.63" reactiontime="+72" points="569">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.79" />
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                    <SPLIT distance="75" swimtime="00:00:44.99" />
                    <SPLIT distance="100" swimtime="00:01:00.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="33" lane="6" heat="1" heatid="10043" swimtime="00:02:13.65" reactiontime="+72" points="562">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.02" />
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="75" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:02.26" />
                    <SPLIT distance="125" swimtime="00:01:19.88" />
                    <SPLIT distance="150" swimtime="00:01:37.66" />
                    <SPLIT distance="175" swimtime="00:01:56.03" />
                    <SPLIT distance="200" swimtime="00:02:13.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Solomon Islands" shortname="SOL" code="SOL" nation="SOL" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="159281" lastname="IRO" firstname="Edgar Richardson" gender="M" birthdate="2000-11-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.90" eventid="14" heat="2" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.52" eventid="31" heat="3" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="80" lane="2" heat="2" heatid="20014" swimtime="00:00:58.43" reactiontime="+65" points="451">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="75" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:00:58.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="71" lane="3" heat="3" heatid="30031" swimtime="00:00:26.62" reactiontime="+66" points="434">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Serbia" shortname="SRB" code="SRB" nation="SRB" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="101098" lastname="STJEPANOVIC" firstname="Velimir" gender="M" birthdate="1993-08-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.43" eventid="14" heat="8" lane="3">
                  <MEETINFO date="2021-09-29" />
                </ENTRY>
                <ENTRY entrytime="00:01:43.30" eventid="44" heat="6" lane="1">
                  <MEETINFO date="2021-09-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="43" lane="3" heat="8" heatid="80014" swimtime="00:00:48.42" reactiontime="+61" points="794">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.26" />
                    <SPLIT distance="50" swimtime="00:00:23.26" />
                    <SPLIT distance="75" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:00:48.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="21" lane="1" heat="6" heatid="60044" swimtime="00:01:44.73" reactiontime="+64" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.46" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:00:50.99" />
                    <SPLIT distance="125" swimtime="00:01:04.40" />
                    <SPLIT distance="150" swimtime="00:01:17.86" />
                    <SPLIT distance="175" swimtime="00:01:31.32" />
                    <SPLIT distance="200" swimtime="00:01:44.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123413" lastname="CREVAR" firstname="Anja" gender="F" birthdate="2000-05-24">
              <ENTRIES>
                <ENTRY entrytime="00:02:12.28" eventid="20" heat="4" lane="1">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:04:09.05" eventid="1" heat="2" lane="6">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
                <ENTRY entrytime="00:04:40.13" eventid="36" heat="2" lane="5">
                  <MEETINFO date="2021-10-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="21" lane="1" heat="4" heatid="40020" swimtime="00:02:12.43" reactiontime="+66" points="736">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="75" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:02.65" />
                    <SPLIT distance="125" swimtime="00:01:19.84" />
                    <SPLIT distance="150" swimtime="00:01:36.99" />
                    <SPLIT distance="175" swimtime="00:01:54.74" />
                    <SPLIT distance="200" swimtime="00:02:12.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="15" lane="6" heat="2" heatid="20001" swimtime="00:04:08.62" reactiontime="+65" points="832">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="75" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:00:59.93" />
                    <SPLIT distance="125" swimtime="00:01:15.55" />
                    <SPLIT distance="150" swimtime="00:01:31.11" />
                    <SPLIT distance="175" swimtime="00:01:46.97" />
                    <SPLIT distance="200" swimtime="00:02:02.80" />
                    <SPLIT distance="225" swimtime="00:02:18.65" />
                    <SPLIT distance="250" swimtime="00:02:34.26" />
                    <SPLIT distance="275" swimtime="00:02:49.99" />
                    <SPLIT distance="300" swimtime="00:03:05.70" />
                    <SPLIT distance="325" swimtime="00:03:21.55" />
                    <SPLIT distance="350" swimtime="00:03:37.38" />
                    <SPLIT distance="375" swimtime="00:03:53.45" />
                    <SPLIT distance="400" swimtime="00:04:08.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="-1" lane="5" heat="2" heatid="20036" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Sri Lanka" shortname="SRI" code="SRI" nation="SRI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="108959" lastname="JASINGHE" firstname="Kiran" gender="M" birthdate="1997-07-13">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.81" eventid="16" heat="3" lane="3">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:56.33" eventid="23" heat="2" lane="7">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="49" lane="3" heat="3" heatid="30016" swimtime="00:01:01.60" reactiontime="+61" points="722">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="75" swimtime="00:00:45.16" />
                    <SPLIT distance="100" swimtime="00:01:01.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="32" lane="7" heat="2" heatid="20023" swimtime="00:00:56.61" reactiontime="+58" points="659">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:26.08" />
                    <SPLIT distance="75" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:00:56.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124808" lastname="PEIRIS" firstname="Dimuth Akalanka" gender="M" birthdate="2000-01-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:25.31" eventid="19" heat="2" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.89" eventid="5" heat="4" lane="7">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="-1" lane="3" heat="2" heatid="20019" swimtime="NT" status="DNS" />
                <RESULT eventid="5" place="-1" lane="7" heat="4" heatid="40005" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="166330" lastname="SENAVIRATHNE" firstname="Ganga" gender="F" birthdate="2003-05-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.51" eventid="2" heat="2" lane="1">
                  <MEETINFO date="2022-10-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.92" eventid="18" heat="3" lane="8">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="-1" lane="1" heat="2" heatid="20002" swimtime="NT" status="DNS" />
                <RESULT eventid="18" place="-1" lane="8" heat="3" heatid="30018" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="149504" lastname="SAMARAKOON" firstname="Ramudi" gender="F" birthdate="2002-11-12">
              <ENTRIES>
                <ENTRY entrytime="00:01:14.54" eventid="15" heat="2" lane="4">
                  <MEETINFO date="2022-10-07" />
                </ENTRY>
                <ENTRY entrytime="00:02:45.53" eventid="28" heat="1" lane="2">
                  <MEETINFO date="2022-10-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="-1" lane="4" heat="2" heatid="20015" swimtime="NT" status="DNS" />
                <RESULT eventid="28" place="-1" lane="2" heat="1" heatid="10028" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Sudan" shortname="SUD" code="SUD" nation="SUD" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="130583" lastname="ABASS" firstname="Abobakr" gender="M" birthdate="1998-11-01">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="3" heat="1" lane="3" />
                <ENTRY entrytime="00:00:28.51" eventid="41" heat="4" lane="8">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="-1" lane="3" heat="1" heatid="10003" swimtime="NT" status="DNS" />
                <RESULT eventid="41" place="46" lane="8" heat="4" heatid="40041" swimtime="00:00:28.44" reactiontime="+66" points="675">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196954" lastname="SALEEM" firstname="Ziyad" gender="M" birthdate="2003-03-24">
              <ENTRIES>
                <ENTRY entrytime="00:02:01.05" eventid="46" heat="1" lane="5">
                  <MEETINFO date="2022-06-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.30" eventid="19" heat="2" lane="5">
                  <MEETINFO date="2021-10-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="-1" lane="5" heat="1" heatid="10046" swimtime="NT" status="DNS" />
                <RESULT eventid="19" place="-1" lane="5" heat="2" heatid="20019" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Switzerland" shortname="SUI" code="SUI" nation="SUI" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="157496" lastname="BOLLIN" firstname="Thierry" gender="M" birthdate="2000-01-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.31" eventid="3" heat="3" lane="4">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.01" eventid="19" heat="4" lane="8">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="4" lane="4" heat="3" heatid="30003" swimtime="00:00:50.10" reactiontime="+60" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.64" />
                    <SPLIT distance="50" swimtime="00:00:24.21" />
                    <SPLIT distance="75" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="10" lane="5" heat="1" heatid="10203" swimtime="00:00:50.33" reactiontime="+60" points="885">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:24.35" />
                    <SPLIT distance="75" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:00:50.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="17" lane="8" heat="4" heatid="40019" swimtime="00:00:23.48" reactiontime="+61" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:23.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="196736" lastname="PONTI" firstname="Noè" gender="M" birthdate="2001-06-01">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.38" eventid="39" heat="6" lane="4">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:49.81" eventid="21" heat="2" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.52" eventid="5" heat="9" lane="2">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="139" place="4" lane="3" heat="1" heatid="10139" swimtime="00:00:49.25" reactiontime="+69" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.46" />
                    <SPLIT distance="50" swimtime="00:00:22.59" />
                    <SPLIT distance="75" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:00:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="1" lane="4" heat="6" heatid="60039" swimtime="00:00:48.81" reactiontime="+70" points="938">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.66" />
                    <SPLIT distance="50" swimtime="00:00:23.13" />
                    <SPLIT distance="75" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:00:48.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="239" place="2" lane="4" heat="2" heatid="20239" swimtime="00:00:49.07" reactiontime="+66" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.03" />
                    <SPLIT distance="75" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="121" place="3" lane="2" heat="1" heatid="10121" swimtime="00:01:49.42" reactiontime="+67" points="967">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.00" />
                    <SPLIT distance="50" swimtime="00:00:24.41" />
                    <SPLIT distance="75" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:00:52.43" />
                    <SPLIT distance="125" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:20.71" />
                    <SPLIT distance="175" swimtime="00:01:34.89" />
                    <SPLIT distance="200" swimtime="00:01:49.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="5" lane="5" heat="2" heatid="20021" swimtime="00:01:50.69" reactiontime="+66" points="935">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.22" />
                    <SPLIT distance="50" swimtime="00:00:25.08" />
                    <SPLIT distance="75" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:00:53.96" />
                    <SPLIT distance="125" swimtime="00:01:07.94" />
                    <SPLIT distance="150" swimtime="00:01:22.29" />
                    <SPLIT distance="175" swimtime="00:01:36.72" />
                    <SPLIT distance="200" swimtime="00:01:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="105" place="2" lane="3" heat="1" heatid="10105" swimtime="00:00:21.96" reactiontime="+64" points="971">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.04" />
                    <SPLIT distance="50" swimtime="00:00:21.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="1" lane="2" heat="9" heatid="90005" swimtime="00:00:22.01" reactiontime="+66" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.16" />
                    <SPLIT distance="50" swimtime="00:00:22.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="3" lane="4" heat="2" heatid="20205" swimtime="00:00:22.04" reactiontime="+64" points="961">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.14" />
                    <SPLIT distance="50" swimtime="00:00:22.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="161939" lastname="DJAKOVIC" firstname="Antonio" gender="M" birthdate="2002-10-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:42.47" eventid="44" heat="5" lane="6">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:03:36.83" eventid="24" heat="4" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="10" lane="6" heat="5" heatid="50044" swimtime="00:01:43.04" reactiontime="+65" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.14" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                    <SPLIT distance="75" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:00:49.73" />
                    <SPLIT distance="125" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:16.43" />
                    <SPLIT distance="175" swimtime="00:01:29.90" />
                    <SPLIT distance="200" swimtime="00:01:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="124" place="5" lane="7" heat="1" heatid="10124" swimtime="00:03:37.86" reactiontime="+70" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.38" />
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                    <SPLIT distance="75" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:00:52.25" />
                    <SPLIT distance="125" swimtime="00:01:06.05" />
                    <SPLIT distance="150" swimtime="00:01:20.02" />
                    <SPLIT distance="175" swimtime="00:01:34.07" />
                    <SPLIT distance="200" swimtime="00:01:48.11" />
                    <SPLIT distance="225" swimtime="00:02:02.08" />
                    <SPLIT distance="250" swimtime="00:02:16.10" />
                    <SPLIT distance="275" swimtime="00:02:30.16" />
                    <SPLIT distance="300" swimtime="00:02:44.28" />
                    <SPLIT distance="325" swimtime="00:02:58.12" />
                    <SPLIT distance="350" swimtime="00:03:11.96" />
                    <SPLIT distance="375" swimtime="00:03:25.31" />
                    <SPLIT distance="400" swimtime="00:03:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="6" lane="5" heat="4" heatid="40024" swimtime="00:03:38.57" reactiontime="+68" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:00:52.82" />
                    <SPLIT distance="125" swimtime="00:01:06.81" />
                    <SPLIT distance="150" swimtime="00:01:20.76" />
                    <SPLIT distance="175" swimtime="00:01:34.87" />
                    <SPLIT distance="200" swimtime="00:01:48.87" />
                    <SPLIT distance="225" swimtime="00:02:02.90" />
                    <SPLIT distance="250" swimtime="00:02:16.85" />
                    <SPLIT distance="275" swimtime="00:02:30.91" />
                    <SPLIT distance="300" swimtime="00:02:44.73" />
                    <SPLIT distance="325" swimtime="00:02:58.69" />
                    <SPLIT distance="350" swimtime="00:03:12.66" />
                    <SPLIT distance="375" swimtime="00:03:26.26" />
                    <SPLIT distance="400" swimtime="00:03:38.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110668" lastname="MAMIE" firstname="Lisa" gender="F" birthdate="1998-10-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.54" eventid="15" heat="5" lane="8">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:23.27" eventid="28" heat="4" lane="8">
                  <MEETINFO date="2022-08-15" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.75" eventid="40" heat="5" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="21" lane="8" heat="5" heatid="50015" swimtime="00:01:05.56" reactiontime="+70" points="860">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                    <SPLIT distance="75" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:05.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="9" lane="8" heat="4" heatid="40028" swimtime="00:02:20.45" reactiontime="+75" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.74" />
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                    <SPLIT distance="75" swimtime="00:00:49.50" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="125" swimtime="00:01:25.37" />
                    <SPLIT distance="150" swimtime="00:01:43.54" />
                    <SPLIT distance="175" swimtime="00:02:02.01" />
                    <SPLIT distance="200" swimtime="00:02:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="24" lane="8" heat="5" heatid="50040" swimtime="00:00:30.84" reactiontime="+69" points="794">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.17" />
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Slovakia" shortname="SVK" code="SVK" nation="SVK" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="125133" lastname="HALAS" firstname="Adam" gender="M" birthdate="1998-08-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.09" eventid="16" heat="4" lane="5">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.43" eventid="39" heat="5" lane="7">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.26" eventid="41" heat="5" lane="4">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.10" eventid="5" heat="7" lane="2">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:53.20" eventid="23" heat="5" lane="1">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="32" lane="5" heat="4" heatid="40016" swimtime="00:00:59.12" reactiontime="+68" points="817">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                    <SPLIT distance="50" swimtime="00:00:27.49" />
                    <SPLIT distance="75" swimtime="00:00:43.16" />
                    <SPLIT distance="100" swimtime="00:00:59.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="22" lane="7" heat="5" heatid="50039" swimtime="00:00:51.34" reactiontime="+68" points="806">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.04" />
                    <SPLIT distance="50" swimtime="00:00:24.14" />
                    <SPLIT distance="75" swimtime="00:00:37.61" />
                    <SPLIT distance="100" swimtime="00:00:51.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="29" lane="4" heat="5" heatid="50041" swimtime="00:00:27.12" reactiontime="+67" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.42" />
                    <SPLIT distance="50" swimtime="00:00:27.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="37" lane="2" heat="7" heatid="70005" swimtime="00:00:23.29" reactiontime="+66" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="22" lane="1" heat="5" heatid="50023" swimtime="00:00:53.43" reactiontime="+69" points="784">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.69" />
                    <SPLIT distance="50" swimtime="00:00:24.28" />
                    <SPLIT distance="75" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:00:53.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154849" lastname="DUSA" firstname="Matej" gender="M" birthdate="2000-07-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.77" eventid="14" heat="6" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.38" eventid="31" heat="10" lane="8">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="35" lane="3" heat="6" heatid="60014" swimtime="00:00:47.75" reactiontime="+59" points="828">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.40" />
                    <SPLIT distance="50" swimtime="00:00:22.37" />
                    <SPLIT distance="75" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:00:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="16" lane="8" heat="10" heatid="100031" swimtime="00:00:21.29" reactiontime="+60" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:21.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="15" lane="8" heat="2" heatid="20231" swimtime="00:00:21.35" reactiontime="+58" points="841">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.04" />
                    <SPLIT distance="50" swimtime="00:00:21.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101620" lastname="KLOBUCNIK" firstname="Tomas" gender="M" birthdate="1990-06-21">
              <ENTRIES>
                <ENTRY entrytime="00:02:06.45" eventid="29" heat="3" lane="7">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="29" place="-1" lane="7" heat="3" heatid="30029" swimtime="00:02:07.87" status="DSQ" reactiontime="+71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102223" lastname="NAGY" firstname="Richard" gender="M" birthdate="1993-03-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:56.93" eventid="21" heat="2" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:59.28" eventid="7" heat="2" lane="3">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:04:10.32" eventid="37" heat="3" lane="8">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="21" place="17" lane="1" heat="2" heatid="20021" swimtime="00:01:54.92" reactiontime="+70" points="835">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                    <SPLIT distance="75" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:00:54.67" />
                    <SPLIT distance="125" swimtime="00:01:09.40" />
                    <SPLIT distance="150" swimtime="00:01:24.41" />
                    <SPLIT distance="175" swimtime="00:01:39.63" />
                    <SPLIT distance="200" swimtime="00:01:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="20" lane="3" heat="2" heatid="20007" swimtime="00:01:57.13" reactiontime="+69" points="819">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                    <SPLIT distance="75" swimtime="00:00:41.26" />
                    <SPLIT distance="100" swimtime="00:00:55.88" />
                    <SPLIT distance="125" swimtime="00:01:12.81" />
                    <SPLIT distance="150" swimtime="00:01:29.62" />
                    <SPLIT distance="175" swimtime="00:01:44.11" />
                    <SPLIT distance="200" swimtime="00:01:57.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="8" lane="8" heat="1" heatid="10137" swimtime="00:04:05.57" reactiontime="+73" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:25.79" />
                    <SPLIT distance="75" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:00:55.18" />
                    <SPLIT distance="125" swimtime="00:01:11.56" />
                    <SPLIT distance="150" swimtime="00:01:27.02" />
                    <SPLIT distance="175" swimtime="00:01:42.71" />
                    <SPLIT distance="200" swimtime="00:01:58.16" />
                    <SPLIT distance="225" swimtime="00:02:15.21" />
                    <SPLIT distance="250" swimtime="00:02:32.62" />
                    <SPLIT distance="275" swimtime="00:02:50.35" />
                    <SPLIT distance="300" swimtime="00:03:08.27" />
                    <SPLIT distance="325" swimtime="00:03:23.53" />
                    <SPLIT distance="350" swimtime="00:03:37.63" />
                    <SPLIT distance="375" swimtime="00:03:51.84" />
                    <SPLIT distance="400" swimtime="00:04:05.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="8" lane="8" heat="3" heatid="30037" swimtime="00:04:06.26" reactiontime="+74" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                    <SPLIT distance="75" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:00:55.01" />
                    <SPLIT distance="125" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:27.22" />
                    <SPLIT distance="175" swimtime="00:01:43.06" />
                    <SPLIT distance="200" swimtime="00:01:58.53" />
                    <SPLIT distance="225" swimtime="00:02:15.82" />
                    <SPLIT distance="250" swimtime="00:02:33.41" />
                    <SPLIT distance="275" swimtime="00:02:51.27" />
                    <SPLIT distance="300" swimtime="00:03:09.44" />
                    <SPLIT distance="325" swimtime="00:03:24.39" />
                    <SPLIT distance="350" swimtime="00:03:38.41" />
                    <SPLIT distance="375" swimtime="00:03:52.60" />
                    <SPLIT distance="400" swimtime="00:04:06.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197033" lastname="POLIACIK" firstname="Jakub" gender="M" birthdate="2004-09-21">
              <ENTRIES>
                <ENTRY entrytime="00:01:45.76" eventid="44" heat="3" lane="3">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:03:48.88" eventid="24" heat="2" lane="2">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:07:59.75" eventid="42" heat="1" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="33" lane="3" heat="3" heatid="30044" swimtime="00:01:47.48" reactiontime="+67" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:00:51.00" />
                    <SPLIT distance="125" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:18.85" />
                    <SPLIT distance="175" swimtime="00:01:33.12" />
                    <SPLIT distance="200" swimtime="00:01:47.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="24" lane="2" heat="2" heatid="20024" swimtime="00:03:49.93" reactiontime="+67" points="786">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:38.95" />
                    <SPLIT distance="100" swimtime="00:00:53.09" />
                    <SPLIT distance="125" swimtime="00:01:07.41" />
                    <SPLIT distance="150" swimtime="00:01:21.89" />
                    <SPLIT distance="175" swimtime="00:01:36.56" />
                    <SPLIT distance="200" swimtime="00:01:51.21" />
                    <SPLIT distance="225" swimtime="00:02:06.08" />
                    <SPLIT distance="250" swimtime="00:02:21.21" />
                    <SPLIT distance="275" swimtime="00:02:36.18" />
                    <SPLIT distance="300" swimtime="00:02:51.09" />
                    <SPLIT distance="325" swimtime="00:03:05.87" />
                    <SPLIT distance="350" swimtime="00:03:20.67" />
                    <SPLIT distance="375" swimtime="00:03:35.57" />
                    <SPLIT distance="400" swimtime="00:03:49.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="19" lane="3" heat="1" heatid="10042" swimtime="00:08:05.91" reactiontime="+67" points="759">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.71" />
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                    <SPLIT distance="75" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:00:56.57" />
                    <SPLIT distance="125" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:26.51" />
                    <SPLIT distance="175" swimtime="00:01:41.66" />
                    <SPLIT distance="200" swimtime="00:01:56.87" />
                    <SPLIT distance="225" swimtime="00:02:12.01" />
                    <SPLIT distance="250" swimtime="00:02:27.26" />
                    <SPLIT distance="275" swimtime="00:02:42.53" />
                    <SPLIT distance="300" swimtime="00:02:57.80" />
                    <SPLIT distance="325" swimtime="00:03:13.15" />
                    <SPLIT distance="350" swimtime="00:03:28.65" />
                    <SPLIT distance="375" swimtime="00:03:44.20" />
                    <SPLIT distance="400" swimtime="00:03:59.75" />
                    <SPLIT distance="425" swimtime="00:04:15.20" />
                    <SPLIT distance="450" swimtime="00:04:30.58" />
                    <SPLIT distance="475" swimtime="00:04:46.11" />
                    <SPLIT distance="500" swimtime="00:05:01.60" />
                    <SPLIT distance="525" swimtime="00:05:17.23" />
                    <SPLIT distance="550" swimtime="00:05:32.73" />
                    <SPLIT distance="575" swimtime="00:05:48.35" />
                    <SPLIT distance="600" swimtime="00:06:03.80" />
                    <SPLIT distance="625" swimtime="00:06:19.11" />
                    <SPLIT distance="650" swimtime="00:06:34.40" />
                    <SPLIT distance="675" swimtime="00:06:49.62" />
                    <SPLIT distance="700" swimtime="00:07:05.11" />
                    <SPLIT distance="725" swimtime="00:07:20.54" />
                    <SPLIT distance="750" swimtime="00:07:35.84" />
                    <SPLIT distance="775" swimtime="00:07:51.26" />
                    <SPLIT distance="800" swimtime="00:08:05.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110770" lastname="PODMANIKOVA" firstname="Andrea" gender="F" birthdate="1998-02-23">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.25" eventid="15" heat="5" lane="7">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:21.15" eventid="28" heat="5" lane="2">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:29.89" eventid="40" heat="5" lane="6">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="18" lane="7" heat="5" heatid="50015" swimtime="00:01:05.31" reactiontime="+69" points="870">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.14" />
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="75" swimtime="00:00:48.06" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="20" lane="2" heat="5" heatid="50028" swimtime="00:02:24.12" reactiontime="+75" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.57" />
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="75" swimtime="00:00:49.37" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="125" swimtime="00:01:25.84" />
                    <SPLIT distance="150" swimtime="00:01:44.57" />
                    <SPLIT distance="175" swimtime="00:02:03.97" />
                    <SPLIT distance="200" swimtime="00:02:24.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="14" lane="6" heat="5" heatid="50040" swimtime="00:00:30.14" reactiontime="+67" points="850">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="15" lane="1" heat="1" heatid="10240" swimtime="00:00:30.21" reactiontime="+68" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156377" lastname="RIPKOVÁ" firstname="Zora" gender="F" birthdate="2002-07-14">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.09" eventid="38" heat="1" lane="6">
                  <MEETINFO date="2022-03-31" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.41" eventid="20" heat="3" lane="7">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="23" lane="6" heat="1" heatid="10038" swimtime="00:00:59.39" reactiontime="+69" points="776">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.02" />
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                    <SPLIT distance="75" swimtime="00:00:43.07" />
                    <SPLIT distance="100" swimtime="00:00:59.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="19" lane="7" heat="3" heatid="30020" swimtime="00:02:11.72" reactiontime="+70" points="748">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                    <SPLIT distance="75" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="125" swimtime="00:01:19.11" />
                    <SPLIT distance="150" swimtime="00:01:36.39" />
                    <SPLIT distance="175" swimtime="00:01:53.79" />
                    <SPLIT distance="200" swimtime="00:02:11.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="198066" lastname="IVANOVA" firstname="Teresa" gender="F" birthdate="2003-09-19">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:54.97" eventid="13" heat="6" lane="3">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:29.02" eventid="18" heat="4" lane="8">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="27" lane="3" heat="6" heatid="60013" swimtime="00:00:54.42" reactiontime="+71" points="787">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.31" />
                    <SPLIT distance="50" swimtime="00:00:25.92" />
                    <SPLIT distance="75" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:00:54.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="33" lane="8" heat="4" heatid="40018" swimtime="00:00:28.29" reactiontime="+67" points="712">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150563" lastname="POTOCKÁ" firstname="Tamara" gender="F" birthdate="2002-08-15">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.33" eventid="45" heat="4" lane="8">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:01:00.52" eventid="22" heat="2" lane="2">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="45" place="25" lane="8" heat="4" heatid="40045" swimtime="00:02:08.61" reactiontime="+60" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.15" />
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="75" swimtime="00:00:46.05" />
                    <SPLIT distance="100" swimtime="00:01:02.60" />
                    <SPLIT distance="125" swimtime="00:01:19.02" />
                    <SPLIT distance="150" swimtime="00:01:35.56" />
                    <SPLIT distance="175" swimtime="00:01:52.19" />
                    <SPLIT distance="200" swimtime="00:02:08.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="13" lane="2" heat="2" heatid="20022" swimtime="00:00:59.69" reactiontime="+70" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.29" />
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                    <SPLIT distance="75" swimtime="00:00:44.99" />
                    <SPLIT distance="100" swimtime="00:00:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="13" lane="1" heat="2" heatid="20222" swimtime="00:00:59.55" reactiontime="+69" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.27" />
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="75" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:00:59.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150565" lastname="TRNÍKOVÁ" firstname="Nikoleta" gender="F" birthdate="2002-07-29">
              <ENTRIES>
                <ENTRY entrytime="00:02:23.04" eventid="28" heat="3" lane="1">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:11.41" eventid="6" heat="4" lane="8">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:04:37.69" eventid="36" heat="3" lane="8">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="21" lane="1" heat="3" heatid="30028" swimtime="00:02:24.62" reactiontime="+63" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.88" />
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="75" swimtime="00:00:50.78" />
                    <SPLIT distance="100" swimtime="00:01:09.18" />
                    <SPLIT distance="125" swimtime="00:01:27.80" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                    <SPLIT distance="175" swimtime="00:02:05.44" />
                    <SPLIT distance="200" swimtime="00:02:24.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="27" lane="8" heat="4" heatid="40006" swimtime="00:02:13.00" reactiontime="+64" points="769">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="75" swimtime="00:00:47.22" />
                    <SPLIT distance="100" swimtime="00:01:03.92" />
                    <SPLIT distance="125" swimtime="00:01:22.59" />
                    <SPLIT distance="150" swimtime="00:01:41.30" />
                    <SPLIT distance="175" swimtime="00:01:57.95" />
                    <SPLIT distance="200" swimtime="00:02:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="15" lane="8" heat="3" heatid="30036" swimtime="00:04:40.09" reactiontime="+65" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="75" swimtime="00:00:47.79" />
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="125" swimtime="00:01:24.14" />
                    <SPLIT distance="150" swimtime="00:01:41.62" />
                    <SPLIT distance="175" swimtime="00:01:59.47" />
                    <SPLIT distance="200" swimtime="00:02:17.00" />
                    <SPLIT distance="225" swimtime="00:02:36.46" />
                    <SPLIT distance="250" swimtime="00:02:55.63" />
                    <SPLIT distance="275" swimtime="00:03:14.92" />
                    <SPLIT distance="300" swimtime="00:03:34.45" />
                    <SPLIT distance="325" swimtime="00:03:51.47" />
                    <SPLIT distance="350" swimtime="00:04:07.73" />
                    <SPLIT distance="375" swimtime="00:04:24.18" />
                    <SPLIT distance="400" swimtime="00:04:40.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156376" lastname="CIBULKOVÁ" firstname="Martina" gender="F" birthdate="2003-11-10">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.48" eventid="43" heat="2" lane="5">
                  <MEETINFO date="2022-10-15" />
                </ENTRY>
                <ENTRY entrytime="00:04:22.80" eventid="1" heat="1" lane="5">
                  <MEETINFO date="2022-11-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="24" lane="5" heat="2" heatid="20043" swimtime="00:02:02.20" reactiontime="+70" points="735">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="75" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:00:58.23" />
                    <SPLIT distance="125" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:29.52" />
                    <SPLIT distance="175" swimtime="00:01:45.87" />
                    <SPLIT distance="200" swimtime="00:02:02.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="23" lane="5" heat="1" heatid="10001" swimtime="00:04:19.76" reactiontime="+69" points="730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="75" swimtime="00:00:44.24" />
                    <SPLIT distance="100" swimtime="00:01:00.13" />
                    <SPLIT distance="125" swimtime="00:01:16.09" />
                    <SPLIT distance="150" swimtime="00:01:32.54" />
                    <SPLIT distance="175" swimtime="00:01:48.77" />
                    <SPLIT distance="200" swimtime="00:02:05.41" />
                    <SPLIT distance="225" swimtime="00:02:21.72" />
                    <SPLIT distance="250" swimtime="00:02:38.50" />
                    <SPLIT distance="275" swimtime="00:02:55.52" />
                    <SPLIT distance="300" swimtime="00:03:12.46" />
                    <SPLIT distance="325" swimtime="00:03:29.42" />
                    <SPLIT distance="350" swimtime="00:03:46.40" />
                    <SPLIT distance="375" swimtime="00:04:03.32" />
                    <SPLIT distance="400" swimtime="00:04:19.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197037" lastname="SLUSNA" firstname="Lillian" gender="F" birthdate="2005-10-27">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:26.54" eventid="4" heat="5" lane="8">
                  <MEETINFO date="2022-10-15" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.77" eventid="30" heat="6" lane="7">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="23" lane="8" heat="5" heatid="50004" swimtime="00:00:26.30" reactiontime="+71" points="796">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.05" />
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="20" lane="7" heat="6" heatid="60030" swimtime="00:00:24.93" reactiontime="+67" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:24.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Slovakia">
              <RESULTS>
                <RESULT eventid="27" place="10" lane="3" heat="3" swimtime="00:01:32.38" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.28" />
                    <SPLIT distance="50" swimtime="00:00:21.58" />
                    <SPLIT distance="75" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:00:43.47" />
                    <SPLIT distance="125" swimtime="00:00:55.18" />
                    <SPLIT distance="150" swimtime="00:01:07.73" />
                    <SPLIT distance="175" swimtime="00:01:19.49" />
                    <SPLIT distance="200" swimtime="00:01:32.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154849" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="125133" reactiontime="+40" />
                    <RELAYPOSITION number="3" athleteid="198066" reactiontime="+46" />
                    <RELAYPOSITION number="4" athleteid="197037" reactiontime="+42" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Slovakia">
              <RESULTS>
                <RESULT eventid="8" place="10" lane="7" heat="2" swimtime="00:03:39.23" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                    <SPLIT distance="75" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:00:55.34" />
                    <SPLIT distance="125" swimtime="00:01:07.55" />
                    <SPLIT distance="150" swimtime="00:01:21.55" />
                    <SPLIT distance="175" swimtime="00:01:35.69" />
                    <SPLIT distance="200" swimtime="00:01:49.80" />
                    <SPLIT distance="225" swimtime="00:02:02.78" />
                    <SPLIT distance="250" swimtime="00:02:16.92" />
                    <SPLIT distance="275" swimtime="00:02:31.19" />
                    <SPLIT distance="300" swimtime="00:02:45.42" />
                    <SPLIT distance="325" swimtime="00:02:57.19" />
                    <SPLIT distance="350" swimtime="00:03:10.91" />
                    <SPLIT distance="375" swimtime="00:03:24.95" />
                    <SPLIT distance="400" swimtime="00:03:39.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197037" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="150563" reactiontime="+42" />
                    <RELAYPOSITION number="3" athleteid="156377" reactiontime="+50" />
                    <RELAYPOSITION number="4" athleteid="198066" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Slovakia">
              <RESULTS>
                <RESULT eventid="47" place="11" lane="8" heat="1" swimtime="00:03:59.50" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="75" swimtime="00:00:43.42" />
                    <SPLIT distance="100" swimtime="00:00:58.73" />
                    <SPLIT distance="125" swimtime="00:01:12.74" />
                    <SPLIT distance="150" swimtime="00:01:29.89" />
                    <SPLIT distance="175" swimtime="00:01:47.59" />
                    <SPLIT distance="200" swimtime="00:02:05.86" />
                    <SPLIT distance="225" swimtime="00:02:18.58" />
                    <SPLIT distance="250" swimtime="00:02:33.44" />
                    <SPLIT distance="275" swimtime="00:02:48.80" />
                    <SPLIT distance="300" swimtime="00:03:05.10" />
                    <SPLIT distance="325" swimtime="00:03:17.00" />
                    <SPLIT distance="350" swimtime="00:03:30.76" />
                    <SPLIT distance="375" swimtime="00:03:45.09" />
                    <SPLIT distance="400" swimtime="00:03:59.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150563" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="110770" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="156377" reactiontime="+31" />
                    <RELAYPOSITION number="4" athleteid="198066" reactiontime="+19" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Slovakia">
              <RESULTS>
                <RESULT eventid="17" place="9" lane="7" heat="2" swimtime="00:08:01.71" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.40" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="75" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:00:58.07" />
                    <SPLIT distance="125" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:28.56" />
                    <SPLIT distance="175" swimtime="00:01:44.35" />
                    <SPLIT distance="200" swimtime="00:01:59.78" />
                    <SPLIT distance="225" swimtime="00:02:12.42" />
                    <SPLIT distance="250" swimtime="00:02:27.09" />
                    <SPLIT distance="275" swimtime="00:02:42.08" />
                    <SPLIT distance="300" swimtime="00:02:57.42" />
                    <SPLIT distance="325" swimtime="00:03:12.41" />
                    <SPLIT distance="350" swimtime="00:03:27.94" />
                    <SPLIT distance="375" swimtime="00:03:43.41" />
                    <SPLIT distance="400" swimtime="00:03:58.46" />
                    <SPLIT distance="425" swimtime="00:04:11.11" />
                    <SPLIT distance="450" swimtime="00:04:26.08" />
                    <SPLIT distance="475" swimtime="00:04:40.96" />
                    <SPLIT distance="500" swimtime="00:04:56.59" />
                    <SPLIT distance="525" swimtime="00:05:12.49" />
                    <SPLIT distance="550" swimtime="00:05:28.91" />
                    <SPLIT distance="575" swimtime="00:05:45.49" />
                    <SPLIT distance="600" swimtime="00:06:01.52" />
                    <SPLIT distance="625" swimtime="00:06:14.73" />
                    <SPLIT distance="650" swimtime="00:06:29.48" />
                    <SPLIT distance="675" swimtime="00:06:44.46" />
                    <SPLIT distance="700" swimtime="00:07:00.00" />
                    <SPLIT distance="725" swimtime="00:07:15.15" />
                    <SPLIT distance="750" swimtime="00:07:30.90" />
                    <SPLIT distance="775" swimtime="00:07:46.39" />
                    <SPLIT distance="800" swimtime="00:08:01.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="156377" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="150563" reactiontime="+42" />
                    <RELAYPOSITION number="3" athleteid="198066" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="156376" reactiontime="+53" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Slovakia">
              <RESULTS>
                <RESULT eventid="25" place="10" lane="3" heat="1" swimtime="00:01:40.78" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:24.61" />
                    <SPLIT distance="75" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:00:50.48" />
                    <SPLIT distance="125" swimtime="00:01:02.74" />
                    <SPLIT distance="150" swimtime="00:01:15.99" />
                    <SPLIT distance="175" swimtime="00:01:27.82" />
                    <SPLIT distance="200" swimtime="00:01:40.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="198066" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="156376" reactiontime="+32" />
                    <RELAYPOSITION number="3" athleteid="156377" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="197037" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Slovakia">
              <RESULTS>
                <RESULT eventid="34" place="11" lane="2" heat="2" swimtime="00:01:48.51" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="75" swimtime="00:00:41.86" />
                    <SPLIT distance="100" swimtime="00:00:58.16" />
                    <SPLIT distance="125" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:24.28" />
                    <SPLIT distance="175" swimtime="00:01:35.74" />
                    <SPLIT distance="200" swimtime="00:01:48.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150563" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="110770" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="197037" reactiontime="+6" />
                    <RELAYPOSITION number="4" athleteid="198066" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Slovakia">
              <RESULTS>
                <RESULT eventid="11" place="15" lane="6" heat="4" swimtime="00:01:42.23" reactiontime="+55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="75" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:00:58.24" />
                    <SPLIT distance="125" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:21.18" />
                    <SPLIT distance="175" swimtime="00:01:31.07" />
                    <SPLIT distance="200" swimtime="00:01:42.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150563" reactiontime="+55" />
                    <RELAYPOSITION number="2" athleteid="110770" reactiontime="+48" />
                    <RELAYPOSITION number="3" athleteid="125133" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="154849" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Sweden" shortname="SWE" code="SWE" nation="SWE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="113443" lastname="PERSSON" firstname="Erik" gender="M" birthdate="1994-01-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.51" eventid="16" heat="6" lane="2">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.18" eventid="29" heat="3" lane="4">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="20" lane="2" heat="6" heatid="60016" swimtime="00:00:58.05" reactiontime="+66" points="863">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.67" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:00:58.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="129" place="5" lane="7" heat="1" heatid="10129" swimtime="00:02:03.19" reactiontime="+67" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                    <SPLIT distance="75" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:00:59.46" />
                    <SPLIT distance="125" swimtime="00:01:15.22" />
                    <SPLIT distance="150" swimtime="00:01:31.06" />
                    <SPLIT distance="175" swimtime="00:01:47.02" />
                    <SPLIT distance="200" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="6" lane="4" heat="3" heatid="30029" swimtime="00:02:04.01" reactiontime="+71" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="75" swimtime="00:00:44.07" />
                    <SPLIT distance="100" swimtime="00:01:00.00" />
                    <SPLIT distance="125" swimtime="00:01:15.86" />
                    <SPLIT distance="150" swimtime="00:01:31.81" />
                    <SPLIT distance="175" swimtime="00:01:47.90" />
                    <SPLIT distance="200" swimtime="00:02:04.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197878" lastname="HOFF" firstname="Oskar" gender="M" birthdate="1998-12-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.35" eventid="39" heat="5" lane="6">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.95" eventid="5" heat="7" lane="3">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:53.82" eventid="23" heat="4" lane="8">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="21" lane="6" heat="5" heatid="50039" swimtime="00:00:51.28" reactiontime="+65" points="808">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.76" />
                    <SPLIT distance="50" swimtime="00:00:23.55" />
                    <SPLIT distance="75" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="31" lane="3" heat="7" heatid="70005" swimtime="00:00:23.01" reactiontime="+63" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.45" />
                    <SPLIT distance="50" swimtime="00:00:23.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="21" lane="8" heat="4" heatid="40023" swimtime="00:00:53.23" reactiontime="+66" points="793">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.71" />
                    <SPLIT distance="75" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:00:53.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="121284" lastname="ELIASSON" firstname="Isak" gender="M" birthdate="1996-01-22">
              <ENTRIES>
                <ENTRY entrytime="00:00:47.37" eventid="14" heat="8" lane="4">
                  <MEETINFO date="2021-11-27" />
                </ENTRY>
                <ENTRY entrytime="00:01:45.18" eventid="44" heat="5" lane="8">
                  <MEETINFO date="2021-11-26" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.60" eventid="31" heat="8" lane="6">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="34" lane="4" heat="8" heatid="80014" swimtime="00:00:47.73" reactiontime="+68" points="829">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.84" />
                    <SPLIT distance="50" swimtime="00:00:22.98" />
                    <SPLIT distance="75" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="25" lane="8" heat="5" heatid="50044" swimtime="00:01:45.17" reactiontime="+70" points="843">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.35" />
                    <SPLIT distance="50" swimtime="00:00:23.98" />
                    <SPLIT distance="75" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:00:50.20" />
                    <SPLIT distance="125" swimtime="00:01:03.51" />
                    <SPLIT distance="150" swimtime="00:01:17.03" />
                    <SPLIT distance="175" swimtime="00:01:31.00" />
                    <SPLIT distance="200" swimtime="00:01:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="29" lane="6" heat="8" heatid="80031" swimtime="00:00:21.47" reactiontime="+68" points="827">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.37" />
                    <SPLIT distance="50" swimtime="00:00:21.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124194" lastname="JOHANSSON" firstname="Victor" gender="M" birthdate="1998-09-13">
              <ENTRIES>
                <ENTRY entrytime="00:15:05.53" eventid="10" heat="1" lane="5">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
                <ENTRY entrytime="00:03:51.29" eventid="24" heat="2" lane="7">
                  <MEETINFO date="2022-08-17" />
                </ENTRY>
                <ENTRY entrytime="00:07:49.14" eventid="42" heat="2" lane="3">
                  <MEETINFO date="2021-07-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="-1" lane="5" heat="1" heatid="10010" swimtime="NT" status="DNS" />
                <RESULT eventid="24" place="-1" lane="7" heat="2" heatid="20024" swimtime="NT" status="DNS" />
                <RESULT eventid="142" place="-1" lane="3" heat="2" heatid="20042" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100526" lastname="HANSSON" firstname="Louise" gender="F" birthdate="1996-11-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.20" eventid="2" heat="6" lane="4">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.02" eventid="38" heat="3" lane="4">
                  <MEETINFO date="2022-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.83" eventid="18" heat="7" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="00:00:58.12" eventid="22" heat="3" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="5" lane="6" heat="1" heatid="10102" swimtime="00:00:55.89" reactiontime="+60" points="947">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.66" />
                    <SPLIT distance="75" swimtime="00:00:41.20" />
                    <SPLIT distance="100" swimtime="00:00:55.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="1" lane="4" heat="6" heatid="60002" swimtime="00:00:56.04" reactiontime="+62" points="939">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                    <SPLIT distance="75" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:00:56.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="3" lane="4" heat="2" heatid="20202" swimtime="00:00:56.08" reactiontime="+62" points="937">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.95" />
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                    <SPLIT distance="75" swimtime="00:00:41.60" />
                    <SPLIT distance="100" swimtime="00:00:56.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="138" place="3" lane="5" heat="1" heatid="10138" swimtime="00:00:54.87" reactiontime="+71" points="984">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:25.61" />
                    <SPLIT distance="75" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:00:54.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="1" lane="4" heat="3" heatid="30038" swimtime="00:00:55.74" reactiontime="+68" points="939">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                    <SPLIT distance="75" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:00:55.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="2" lane="4" heat="2" heatid="20238" swimtime="00:00:55.78" reactiontime="+69" points="937">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="75" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:00:55.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="5" lane="2" heat="1" heatid="10118" swimtime="00:00:26.00" reactiontime="+61" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.77" />
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="4" lane="5" heat="7" heatid="70018" swimtime="00:00:26.07" reactiontime="+60" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.85" />
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="5" lane="3" heat="1" heatid="10218" swimtime="00:00:25.99" reactiontime="+60" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="122" place="3" lane="5" heat="1" heatid="10122" swimtime="00:00:57.68" reactiontime="+67" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                    <SPLIT distance="75" swimtime="00:00:43.49" />
                    <SPLIT distance="100" swimtime="00:00:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="1" lane="4" heat="3" heatid="30022" swimtime="00:00:57.98" reactiontime="+67" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.67" />
                    <SPLIT distance="50" swimtime="00:00:25.96" />
                    <SPLIT distance="75" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:00:57.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="2" lane="4" heat="2" heatid="20222" swimtime="00:00:58.05" reactiontime="+69" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.57" />
                    <SPLIT distance="50" swimtime="00:00:26.03" />
                    <SPLIT distance="75" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:00:58.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129785" lastname="ROSVALL" firstname="Hanna" gender="F" birthdate="2000-02-10">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.56" eventid="2" heat="5" lane="7">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.82" eventid="45" heat="5" lane="1">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:26.39" eventid="18" heat="6" lane="2">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="4" lane="7" heat="5" heatid="50002" swimtime="00:00:56.57" reactiontime="+59" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                    <SPLIT distance="75" swimtime="00:00:42.00" />
                    <SPLIT distance="100" swimtime="00:00:56.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="9" lane="5" heat="1" heatid="10202" swimtime="00:00:56.59" reactiontime="+59" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                    <SPLIT distance="75" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:00:56.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="10" lane="1" heat="5" heatid="50045" swimtime="00:02:04.37" reactiontime="+59" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.97" />
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="75" swimtime="00:00:45.24" />
                    <SPLIT distance="100" swimtime="00:01:01.30" />
                    <SPLIT distance="125" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:01:33.05" />
                    <SPLIT distance="175" swimtime="00:01:49.04" />
                    <SPLIT distance="200" swimtime="00:02:04.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="6" lane="7" heat="1" heatid="10118" swimtime="00:00:26.05" reactiontime="+58" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="4" lane="2" heat="6" heatid="60018" swimtime="00:00:26.07" reactiontime="+59" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="6" lane="3" heat="2" heatid="20218" swimtime="00:00:26.01" reactiontime="+60" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:26.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124193" lastname="HANSSON" firstname="Sophie" gender="F" birthdate="1998-08-02">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.50" eventid="15" heat="7" lane="5">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:02:18.13" eventid="28" heat="4" lane="4">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:29.55" eventid="40" heat="5" lane="5">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="9" lane="5" heat="7" heatid="70015" swimtime="00:01:04.64" reactiontime="+71" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="75" swimtime="00:00:47.34" />
                    <SPLIT distance="100" swimtime="00:01:04.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="10" lane="2" heat="2" heatid="20215" swimtime="00:01:04.88" reactiontime="+70" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.95" />
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="75" swimtime="00:00:47.69" />
                    <SPLIT distance="100" swimtime="00:01:04.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="-1" lane="4" heat="4" heatid="40028" swimtime="NT" status="DNS" />
                <RESULT eventid="40" place="-1" lane="5" heat="5" heatid="50040" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197607" lastname="THORMALM" firstname="Klara" gender="F" birthdate="1998-03-29">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:05.82" eventid="15" heat="4" lane="5">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:29.96" eventid="40" heat="6" lane="2">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="23" lane="5" heat="4" heatid="40015" swimtime="00:01:05.85" reactiontime="+74" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="75" swimtime="00:00:47.88" />
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="13" lane="2" heat="6" heatid="60040" swimtime="00:00:30.06" reactiontime="+71" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.69" />
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="12" lane="1" heat="2" heatid="20240" swimtime="00:00:30.01" reactiontime="+73" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101062" lastname="COLEMAN" firstname="Michelle" gender="F" birthdate="1993-10-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.94" eventid="13" heat="7" lane="3">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:23.84" eventid="30" heat="7" lane="5">
                  <MEETINFO date="2021-09-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="10" lane="3" heat="7" heatid="70013" swimtime="00:00:52.67" reactiontime="+68" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                    <SPLIT distance="50" swimtime="00:00:25.58" />
                    <SPLIT distance="75" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:00:52.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="10" lane="2" heat="1" heatid="10213" swimtime="00:00:52.44" reactiontime="+68" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                    <SPLIT distance="75" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:00:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="5" lane="3" heat="1" heatid="10130" swimtime="00:00:23.72" reactiontime="+70" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:23.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="7" lane="5" heat="7" heatid="70030" swimtime="00:00:23.94" reactiontime="+69" points="878">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:23.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="3" lane="6" heat="2" heatid="20230" swimtime="00:00:23.77" reactiontime="+67" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:23.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129915" lastname="JUNEVIK" firstname="Sara" gender="F" birthdate="2000-02-14">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.72" eventid="13" heat="7" lane="1">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:25.36" eventid="4" heat="4" lane="6">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="12" lane="1" heat="7" heatid="70013" swimtime="00:00:52.91" reactiontime="+76" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                    <SPLIT distance="75" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:00:52.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="11" lane="7" heat="1" heatid="10213" swimtime="00:00:52.50" reactiontime="+68" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:24.98" />
                    <SPLIT distance="75" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="104" place="8" lane="8" heat="1" heatid="10104" swimtime="00:00:25.18" reactiontime="+71" points="907">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:25.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="3" lane="6" heat="4" heatid="40004" swimtime="00:00:25.04" reactiontime="+71" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.49" />
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="8" lane="5" heat="2" heatid="20204" swimtime="00:00:25.13" reactiontime="+72" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156861" lastname="FAST" firstname="Emelie" gender="F" birthdate="2004-02-20">
              <ENTRIES>
                <ENTRY entrytime="00:02:22.02" eventid="28" heat="4" lane="1">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="00:02:10.82" eventid="6" heat="4" lane="1">
                  <MEETINFO date="2021-11-24" />
                </ENTRY>
                <ENTRY entrytime="00:00:59.50" eventid="22" heat="4" lane="6">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="17" lane="1" heat="4" heatid="40028" swimtime="00:02:22.22" reactiontime="+66" points="847">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.23" />
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="75" swimtime="00:00:49.05" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="125" swimtime="00:01:25.69" />
                    <SPLIT distance="150" swimtime="00:01:44.06" />
                    <SPLIT distance="175" swimtime="00:02:03.11" />
                    <SPLIT distance="200" swimtime="00:02:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="22" lane="1" heat="4" heatid="40006" swimtime="00:02:10.95" reactiontime="+63" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.34" />
                    <SPLIT distance="50" swimtime="00:00:27.61" />
                    <SPLIT distance="75" swimtime="00:00:44.75" />
                    <SPLIT distance="100" swimtime="00:01:01.55" />
                    <SPLIT distance="125" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:01:38.28" />
                    <SPLIT distance="175" swimtime="00:01:55.04" />
                    <SPLIT distance="200" swimtime="00:02:10.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="22" place="12" lane="6" heat="4" heatid="40022" swimtime="00:00:59.53" reactiontime="+64" points="855">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.21" />
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                    <SPLIT distance="75" swimtime="00:00:44.47" />
                    <SPLIT distance="100" swimtime="00:00:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="222" place="14" lane="7" heat="1" heatid="10222" swimtime="00:00:59.61" reactiontime="+67" points="851">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.20" />
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                    <SPLIT distance="75" swimtime="00:00:44.66" />
                    <SPLIT distance="100" swimtime="00:00:59.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197610" lastname="AASTEDT" firstname="Sofia" gender="F" birthdate="2003-11-13">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:58.00" eventid="43" heat="3" lane="1">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="20" lane="1" heat="3" heatid="30043" swimtime="00:01:58.04" reactiontime="+72" points="816">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.01" />
                    <SPLIT distance="50" swimtime="00:00:27.42" />
                    <SPLIT distance="75" swimtime="00:00:42.24" />
                    <SPLIT distance="100" swimtime="00:00:57.30" />
                    <SPLIT distance="125" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:27.72" />
                    <SPLIT distance="175" swimtime="00:01:43.11" />
                    <SPLIT distance="200" swimtime="00:01:58.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Sweden">
              <RESULTS>
                <RESULT eventid="27" place="9" lane="5" heat="2" swimtime="00:01:32.34" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.90" />
                    <SPLIT distance="50" swimtime="00:00:22.46" />
                    <SPLIT distance="75" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:00:43.25" />
                    <SPLIT distance="125" swimtime="00:00:54.86" />
                    <SPLIT distance="150" swimtime="00:01:07.53" />
                    <SPLIT distance="175" swimtime="00:01:19.32" />
                    <SPLIT distance="200" swimtime="00:01:32.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197878" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="121284" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="197610" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="197607" reactiontime="+26" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Sweden">
              <RESULTS>
                <RESULT eventid="108" place="4" lane="7" heat="1" swimtime="00:03:29.35" reactiontime="+71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:24.97" />
                    <SPLIT distance="75" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:00:52.46" />
                    <SPLIT distance="125" swimtime="00:01:03.86" />
                    <SPLIT distance="150" swimtime="00:01:17.01" />
                    <SPLIT distance="175" swimtime="00:01:30.62" />
                    <SPLIT distance="200" swimtime="00:01:44.22" />
                    <SPLIT distance="225" swimtime="00:01:56.09" />
                    <SPLIT distance="250" swimtime="00:02:09.18" />
                    <SPLIT distance="275" swimtime="00:02:22.81" />
                    <SPLIT distance="300" swimtime="00:02:36.37" />
                    <SPLIT distance="325" swimtime="00:02:48.20" />
                    <SPLIT distance="350" swimtime="00:03:01.69" />
                    <SPLIT distance="375" swimtime="00:03:15.56" />
                    <SPLIT distance="400" swimtime="00:03:29.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129915" reactiontime="+71" />
                    <RELAYPOSITION number="2" athleteid="101062" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="100526" reactiontime="+60" />
                    <RELAYPOSITION number="4" athleteid="197610" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="6" lane="5" heat="2" swimtime="00:03:33.17" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.06" />
                    <SPLIT distance="50" swimtime="00:00:25.23" />
                    <SPLIT distance="75" swimtime="00:00:38.88" />
                    <SPLIT distance="100" swimtime="00:00:52.79" />
                    <SPLIT distance="125" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:18.49" />
                    <SPLIT distance="175" swimtime="00:01:32.59" />
                    <SPLIT distance="200" swimtime="00:01:46.44" />
                    <SPLIT distance="225" swimtime="00:01:58.21" />
                    <SPLIT distance="250" swimtime="00:02:12.26" />
                    <SPLIT distance="275" swimtime="00:02:26.74" />
                    <SPLIT distance="300" swimtime="00:02:40.94" />
                    <SPLIT distance="325" swimtime="00:02:52.48" />
                    <SPLIT distance="350" swimtime="00:03:05.68" />
                    <SPLIT distance="375" swimtime="00:03:19.49" />
                    <SPLIT distance="400" swimtime="00:03:33.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129915" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="197610" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="197607" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="101062" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Sweden">
              <RESULTS>
                <RESULT eventid="147" place="5" lane="6" heat="1" swimtime="00:03:47.84" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.24" />
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                    <SPLIT distance="75" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:00:56.37" />
                    <SPLIT distance="125" swimtime="00:01:09.90" />
                    <SPLIT distance="150" swimtime="00:01:26.52" />
                    <SPLIT distance="175" swimtime="00:01:43.67" />
                    <SPLIT distance="200" swimtime="00:02:01.33" />
                    <SPLIT distance="225" swimtime="00:02:12.61" />
                    <SPLIT distance="250" swimtime="00:02:26.37" />
                    <SPLIT distance="275" swimtime="00:02:40.73" />
                    <SPLIT distance="300" swimtime="00:02:55.90" />
                    <SPLIT distance="325" swimtime="00:03:07.19" />
                    <SPLIT distance="350" swimtime="00:03:20.08" />
                    <SPLIT distance="375" swimtime="00:03:33.71" />
                    <SPLIT distance="400" swimtime="00:03:47.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129785" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="124193" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="100526" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="101062" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="4" lane="4" heat="2" swimtime="00:03:52.49" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.11" />
                    <SPLIT distance="50" swimtime="00:00:27.22" />
                    <SPLIT distance="75" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:00:56.84" />
                    <SPLIT distance="125" swimtime="00:01:10.60" />
                    <SPLIT distance="150" swimtime="00:01:27.22" />
                    <SPLIT distance="175" swimtime="00:01:44.51" />
                    <SPLIT distance="200" swimtime="00:02:02.11" />
                    <SPLIT distance="225" swimtime="00:02:13.47" />
                    <SPLIT distance="250" swimtime="00:02:27.82" />
                    <SPLIT distance="275" swimtime="00:02:42.68" />
                    <SPLIT distance="300" swimtime="00:02:58.16" />
                    <SPLIT distance="325" swimtime="00:03:10.36" />
                    <SPLIT distance="350" swimtime="00:03:24.10" />
                    <SPLIT distance="375" swimtime="00:03:38.33" />
                    <SPLIT distance="400" swimtime="00:03:52.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100526" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="197607" reactiontime="+10" />
                    <RELAYPOSITION number="3" athleteid="129915" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="197610" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Sweden">
              <RESULTS>
                <RESULT eventid="125" place="4" lane="1" heat="1" swimtime="00:01:35.68" reactiontime="+69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.13" />
                    <SPLIT distance="75" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:00:47.41" />
                    <SPLIT distance="125" swimtime="00:00:58.81" />
                    <SPLIT distance="150" swimtime="00:01:11.19" />
                    <SPLIT distance="175" swimtime="00:01:22.76" />
                    <SPLIT distance="200" swimtime="00:01:35.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129915" reactiontime="+69" />
                    <RELAYPOSITION number="2" athleteid="101062" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="100526" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="124193" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="7" lane="4" heat="1" swimtime="00:01:37.93" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:24.30" />
                    <SPLIT distance="75" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:00:48.83" />
                    <SPLIT distance="125" swimtime="00:01:00.54" />
                    <SPLIT distance="150" swimtime="00:01:13.35" />
                    <SPLIT distance="175" swimtime="00:01:25.22" />
                    <SPLIT distance="200" swimtime="00:01:37.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129915" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="197610" reactiontime="+30" />
                    <RELAYPOSITION number="3" athleteid="124193" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="129785" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="Sweden">
              <RESULTS>
                <RESULT eventid="134" place="3" lane="5" heat="1" swimtime="00:01:42.43" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.78" />
                    <SPLIT distance="50" swimtime="00:00:25.86" />
                    <SPLIT distance="75" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:00:55.20" />
                    <SPLIT distance="125" swimtime="00:01:05.83" />
                    <SPLIT distance="150" swimtime="00:01:19.26" />
                    <SPLIT distance="175" swimtime="00:01:30.22" />
                    <SPLIT distance="200" swimtime="00:01:42.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="100526" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="197607" reactiontime="+12" />
                    <RELAYPOSITION number="3" athleteid="129915" reactiontime="+5" />
                    <RELAYPOSITION number="4" athleteid="101062" reactiontime="+12" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="2" lane="4" heat="2" swimtime="00:01:44.83" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.18" />
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="75" swimtime="00:00:39.74" />
                    <SPLIT distance="100" swimtime="00:00:55.89" />
                    <SPLIT distance="125" swimtime="00:01:06.69" />
                    <SPLIT distance="150" swimtime="00:01:20.31" />
                    <SPLIT distance="175" swimtime="00:01:31.94" />
                    <SPLIT distance="200" swimtime="00:01:44.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129785" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="197607" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="129915" reactiontime="+9" />
                    <RELAYPOSITION number="4" athleteid="197610" reactiontime="+5" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Sweden">
              <RESULTS>
                <RESULT eventid="11" place="9" lane="5" heat="4" swimtime="00:01:39.26" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="75" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:00:55.80" />
                    <SPLIT distance="125" swimtime="00:01:05.75" />
                    <SPLIT distance="150" swimtime="00:01:18.10" />
                    <SPLIT distance="175" swimtime="00:01:28.05" />
                    <SPLIT distance="200" swimtime="00:01:39.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129785" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="197607" reactiontime="+5" />
                    <RELAYPOSITION number="3" athleteid="197878" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="121284" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Eswatini" shortname="SWZ" code="SWZ" nation="SWZ" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="120198" lastname="DLAMINI" firstname="Simanga" gender="M" birthdate="1997-10-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.46" eventid="39" heat="2" lane="2">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.98" eventid="5" heat="3" lane="8">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="53" lane="2" heat="2" heatid="20039" swimtime="00:01:03.90" reactiontime="+69" points="418">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.56" />
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="75" swimtime="00:00:46.39" />
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="63" lane="8" heat="3" heatid="30005" swimtime="00:00:28.70" reactiontime="+70" points="435">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213598" lastname="JELE" firstname="Cameron" gender="M" birthdate="2006-06-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="41" heat="2" lane="7" />
                <ENTRY entrytime="NT" eventid="31" heat="1" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="56" lane="7" heat="2" heatid="20041" swimtime="00:00:34.95" reactiontime="+68" points="363">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="75" lane="4" heat="1" heatid="10031" swimtime="00:00:28.23" reactiontime="+67" points="364">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197306" lastname="YOUNG" firstname="Raya" gender="F" birthdate="2005-11-20">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="2" heat="1" lane="7" />
                <ENTRY entrytime="NT" eventid="18" heat="1" lane="4" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="47" lane="7" heat="1" heatid="10002" swimtime="00:01:18.68" reactiontime="+65" points="339">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.90" />
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="75" swimtime="00:00:58.71" />
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="50" lane="4" heat="1" heatid="10018" swimtime="00:00:35.86" reactiontime="+65" points="349">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.76" />
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Syrian Arab Rep." shortname="SYR" code="SYR" nation="SYR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="128812" lastname="ABBASS" firstname="Omar" gender="M" birthdate="1999-03-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.99" eventid="14" heat="4" lane="6">
                  <MEETINFO date="2022-06-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.50" eventid="44" heat="2" lane="1">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="51" lane="6" heat="4" heatid="40014" swimtime="00:00:50.01" reactiontime="+67" points="720">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:24.08" />
                    <SPLIT distance="75" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="36" lane="1" heat="2" heatid="20044" swimtime="00:01:48.73" reactiontime="+66" points="763">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.12" />
                    <SPLIT distance="50" swimtime="00:00:25.56" />
                    <SPLIT distance="75" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:00:53.07" />
                    <SPLIT distance="125" swimtime="00:01:06.70" />
                    <SPLIT distance="150" swimtime="00:01:20.67" />
                    <SPLIT distance="175" swimtime="00:01:34.86" />
                    <SPLIT distance="200" swimtime="00:01:48.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101441" lastname="KELZI" firstname="Ayman" gender="M" birthdate="1993-01-07">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="19" heat="1" lane="7" />
                <ENTRY entrytime="00:00:24.64" eventid="5" heat="4" lane="2">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="39" lane="7" heat="1" heatid="10019" swimtime="00:00:27.19" reactiontime="+61" points="545">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.58" />
                    <SPLIT distance="50" swimtime="00:00:27.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="52" lane="2" heat="4" heatid="40005" swimtime="00:00:24.34" reactiontime="+69" points="713">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.23" />
                    <SPLIT distance="50" swimtime="00:00:24.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tanzania" shortname="TAN" code="TAN" nation="TAN" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="141971" lastname="SALIBOKO" firstname="Collins" gender="M" birthdate="2002-04-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.62" eventid="39" heat="3" lane="7">
                  <MEETINFO date="2022-08-22" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.54" eventid="14" heat="3" lane="4">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="43" lane="7" heat="3" heatid="30039" swimtime="00:00:55.85" reactiontime="+56" points="626">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:25.87" />
                    <SPLIT distance="75" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:00:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="62" lane="4" heat="3" heatid="30014" swimtime="00:00:51.50" reactiontime="+58" points="660">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:24.78" />
                    <SPLIT distance="75" swimtime="00:00:38.12" />
                    <SPLIT distance="100" swimtime="00:00:51.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101806" lastname="HILAL" firstname="Hilal" gender="M" birthdate="1994-07-12">
              <ENTRIES>
                <ENTRY entrytime="00:00:29.97" eventid="41" heat="3" lane="8">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.38" eventid="31" heat="4" lane="5">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="53" lane="8" heat="3" heatid="30041" swimtime="00:00:30.23" reactiontime="+59" points="562">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="63" lane="5" heat="4" heatid="40031" swimtime="00:00:24.84" reactiontime="+59" points="534">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:24.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197632" lastname="LATIFF" firstname="Sophia" gender="F" birthdate="2006-12-24">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:01:02.71" eventid="13" heat="3" lane="2">
                  <MEETINFO date="2021-10-11" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.41" eventid="30" heat="3" lane="2">
                  <MEETINFO date="2021-10-15" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="55" lane="2" heat="3" heatid="30013" swimtime="00:01:00.97" reactiontime="+82" points="559">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.04" />
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                    <SPLIT distance="75" swimtime="00:00:45.00" />
                    <SPLIT distance="100" swimtime="00:01:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="41" lane="2" heat="3" heatid="30030" swimtime="00:00:27.63" reactiontime="+70" points="571">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197016" lastname="SAVE" firstname="Ria" gender="F" birthdate="2006-11-20">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:34.69" eventid="18" heat="2" lane="6">
                  <MEETINFO date="2021-10-11" />
                </ENTRY>
                <ENTRY entrytime="00:00:40.65" eventid="40" heat="2" lane="3">
                  <MEETINFO date="2021-10-13" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="44" lane="6" heat="2" heatid="20018" swimtime="00:00:32.90" reactiontime="+57" points="453">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="38" lane="3" heat="2" heatid="20040" swimtime="00:00:38.22" reactiontime="+61" points="417">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="United Republic of Tanzania">
              <RESULTS>
                <RESULT eventid="27" place="22" lane="7" heat="2" swimtime="00:01:44.43" reactiontime="+72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="75" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:00:52.60" />
                    <SPLIT distance="125" swimtime="00:01:06.24" />
                    <SPLIT distance="150" swimtime="00:01:21.09" />
                    <SPLIT distance="175" swimtime="00:01:32.30" />
                    <SPLIT distance="200" swimtime="00:01:44.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197632" reactiontime="+72" />
                    <RELAYPOSITION number="2" athleteid="101806" reactiontime="+73" />
                    <RELAYPOSITION number="3" athleteid="197016" reactiontime="+44" />
                    <RELAYPOSITION number="4" athleteid="141971" reactiontime="+39" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="United Republic of Tanzania">
              <RESULTS>
                <RESULT eventid="11" place="26" lane="7" heat="2" swimtime="00:01:55.82" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="75" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:02.94" />
                    <SPLIT distance="125" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:27.99" />
                    <SPLIT distance="175" swimtime="00:01:41.59" />
                    <SPLIT distance="200" swimtime="00:01:55.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197016" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="101806" reactiontime="+42" />
                    <RELAYPOSITION number="3" athleteid="141971" reactiontime="+48" />
                    <RELAYPOSITION number="4" athleteid="197632" reactiontime="+64" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Tonga" shortname="TGA" code="TGA" nation="TGA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="193830" lastname="UHI" firstname="Alan Koti Lopeti" gender="M" birthdate="2005-10-16">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.94" eventid="3" heat="2" lane="7">
                  <MEETINFO date="2022-07-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.79" eventid="19" heat="1" lane="6">
                  <MEETINFO date="2022-07-31" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="37" lane="7" heat="2" heatid="20003" swimtime="00:00:57.39" reactiontime="+71" points="597">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.02" />
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                    <SPLIT distance="75" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:00:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="38" lane="6" heat="1" heatid="10019" swimtime="00:00:26.84" reactiontime="+68" points="567">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="155060" lastname="OHUAFI" firstname="Finau" gender="M" birthdate="2001-01-25">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.13" eventid="39" heat="3" lane="8">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.77" eventid="14" heat="3" lane="5">
                  <MEETINFO date="2021-10-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="50" lane="8" heat="3" heatid="30039" swimtime="00:00:57.66" reactiontime="+71" points="569">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.31" />
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                    <SPLIT distance="75" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:00:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="67" lane="5" heat="3" heatid="30014" swimtime="00:00:52.91" reactiontime="+67" points="608">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                    <SPLIT distance="75" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:00:52.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102008" lastname="PANUVE" firstname="Charissa" gender="F" birthdate="1994-11-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.95" eventid="13" heat="2" lane="5">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:19.53" eventid="43" heat="1" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="57" lane="5" heat="2" heatid="20013" swimtime="00:01:03.34" reactiontime="+57" points="499">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.39" />
                    <SPLIT distance="50" swimtime="00:00:30.20" />
                    <SPLIT distance="75" swimtime="00:00:46.63" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="34" lane="2" heat="1" heatid="10043" swimtime="00:02:17.97" reactiontime="+57" points="511">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.02" />
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="75" swimtime="00:00:49.03" />
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="125" swimtime="00:01:24.19" />
                    <SPLIT distance="150" swimtime="00:01:42.09" />
                    <SPLIT distance="175" swimtime="00:02:00.23" />
                    <SPLIT distance="200" swimtime="00:02:17.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="135581" lastname="DAY" firstname="Noelani Malia" gender="F" birthdate="2003-04-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.75" eventid="18" heat="2" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:28.14" eventid="30" heat="3" lane="6">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="47" lane="5" heat="2" heatid="20018" swimtime="00:00:33.92" reactiontime="+72" points="413">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="43" lane="6" heat="3" heatid="30030" swimtime="00:00:28.18" reactiontime="+71" points="538">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Thailand" shortname="THA" code="THA" nation="THA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="125335" lastname="WONGCHAROEN" firstname="Navaphat" gender="M" birthdate="1997-03-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:52.98" eventid="39" heat="4" lane="3">
                  <MEETINFO date="2022-05-16" />
                </ENTRY>
                <ENTRY entrytime="00:01:56.55" eventid="21" heat="3" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="32" lane="3" heat="4" heatid="40039" swimtime="00:00:52.19" reactiontime="+54" points="767">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.23" />
                    <SPLIT distance="50" swimtime="00:00:24.49" />
                    <SPLIT distance="75" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:00:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="20" lane="1" heat="3" heatid="30021" swimtime="00:01:56.37" reactiontime="+58" points="804">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.80" />
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                    <SPLIT distance="75" swimtime="00:00:40.58" />
                    <SPLIT distance="100" swimtime="00:00:55.32" />
                    <SPLIT distance="125" swimtime="00:01:10.51" />
                    <SPLIT distance="150" swimtime="00:01:25.85" />
                    <SPLIT distance="175" swimtime="00:01:40.90" />
                    <SPLIT distance="200" swimtime="00:01:56.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202649" lastname="THAMMANANTHACHOTE" firstname="Ratthawit" gender="M" birthdate="2002-09-11">
              <ENTRIES>
                <ENTRY entrytime="00:01:59.04" eventid="46" heat="2" lane="8">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:08:08.52" eventid="42" heat="1" lane="6">
                  <MEETINFO date="2022-04-08" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="46" place="24" lane="8" heat="2" heatid="20046" swimtime="00:02:00.85" reactiontime="+62" points="667">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.96" />
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                    <SPLIT distance="75" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:00:57.93" />
                    <SPLIT distance="125" swimtime="00:01:13.28" />
                    <SPLIT distance="150" swimtime="00:01:29.15" />
                    <SPLIT distance="175" swimtime="00:01:45.08" />
                    <SPLIT distance="200" swimtime="00:02:00.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="17" lane="6" heat="1" heatid="10042" swimtime="00:07:55.24" reactiontime="+76" points="812">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                    <SPLIT distance="75" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:00:56.27" />
                    <SPLIT distance="125" swimtime="00:01:10.97" />
                    <SPLIT distance="150" swimtime="00:01:25.80" />
                    <SPLIT distance="175" swimtime="00:01:40.60" />
                    <SPLIT distance="200" swimtime="00:01:55.48" />
                    <SPLIT distance="225" swimtime="00:02:10.13" />
                    <SPLIT distance="250" swimtime="00:02:25.17" />
                    <SPLIT distance="275" swimtime="00:02:40.01" />
                    <SPLIT distance="300" swimtime="00:02:55.17" />
                    <SPLIT distance="325" swimtime="00:03:09.88" />
                    <SPLIT distance="350" swimtime="00:03:24.84" />
                    <SPLIT distance="375" swimtime="00:03:39.79" />
                    <SPLIT distance="400" swimtime="00:03:55.00" />
                    <SPLIT distance="425" swimtime="00:04:09.94" />
                    <SPLIT distance="450" swimtime="00:04:25.07" />
                    <SPLIT distance="475" swimtime="00:04:40.01" />
                    <SPLIT distance="500" swimtime="00:04:55.28" />
                    <SPLIT distance="525" swimtime="00:05:10.33" />
                    <SPLIT distance="550" swimtime="00:05:25.46" />
                    <SPLIT distance="575" swimtime="00:05:40.41" />
                    <SPLIT distance="600" swimtime="00:05:55.66" />
                    <SPLIT distance="625" swimtime="00:06:10.62" />
                    <SPLIT distance="650" swimtime="00:06:25.74" />
                    <SPLIT distance="675" swimtime="00:06:40.75" />
                    <SPLIT distance="700" swimtime="00:06:55.94" />
                    <SPLIT distance="725" swimtime="00:07:10.97" />
                    <SPLIT distance="750" swimtime="00:07:26.11" />
                    <SPLIT distance="775" swimtime="00:07:41.12" />
                    <SPLIT distance="800" swimtime="00:07:55.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202824" lastname="KAEWSRIYONG" firstname="Dulyawat" gender="M" birthdate="2002-08-13">
              <ENTRIES>
                <ENTRY entrytime="00:02:02.89" eventid="7" heat="2" lane="1">
                  <MEETINFO date="2022-05-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:57.49" eventid="23" heat="2" lane="1">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="31" lane="1" heat="2" heatid="20007" swimtime="00:01:59.85" reactiontime="+65" points="765">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.17" />
                    <SPLIT distance="50" swimtime="00:00:24.71" />
                    <SPLIT distance="75" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:00:55.61" />
                    <SPLIT distance="125" swimtime="00:01:12.91" />
                    <SPLIT distance="150" swimtime="00:01:30.60" />
                    <SPLIT distance="175" swimtime="00:01:45.99" />
                    <SPLIT distance="200" swimtime="00:01:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="31" lane="1" heat="2" heatid="20023" swimtime="00:00:54.81" reactiontime="+67" points="726">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.18" />
                    <SPLIT distance="50" swimtime="00:00:25.52" />
                    <SPLIT distance="75" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:00:54.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123228" lastname="PAWAPOTAKO" firstname="Phiangkhwan" gender="F" birthdate="1996-11-14">
              <ENTRIES>
                <ENTRY entrytime="00:02:27.50" eventid="28" heat="2" lane="8">
                  <MEETINFO date="2021-09-18" />
                </ENTRY>
                <ENTRY entrytime="00:02:14.50" eventid="6" heat="2" lane="1">
                  <MEETINFO date="2021-09-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="26" lane="8" heat="2" heatid="20028" swimtime="00:02:28.50" reactiontime="+67" points="744">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.51" />
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="75" swimtime="00:00:51.54" />
                    <SPLIT distance="100" swimtime="00:01:10.25" />
                    <SPLIT distance="125" swimtime="00:01:29.22" />
                    <SPLIT distance="150" swimtime="00:01:48.77" />
                    <SPLIT distance="175" swimtime="00:02:08.37" />
                    <SPLIT distance="200" swimtime="00:02:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="28" lane="1" heat="2" heatid="20006" swimtime="00:02:13.76" reactiontime="+64" points="756">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.28" />
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="75" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:02.98" />
                    <SPLIT distance="125" swimtime="00:01:21.98" />
                    <SPLIT distance="150" swimtime="00:01:41.46" />
                    <SPLIT distance="175" swimtime="00:01:58.33" />
                    <SPLIT distance="200" swimtime="00:02:13.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="109148" lastname="SRISA - ARD" firstname="Jenjira" gender="F" birthdate="1995-04-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:30.53" eventid="40" heat="7" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.19" eventid="4" heat="5" lane="7">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.78" eventid="30" heat="8" lane="1">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="21" lane="8" heat="7" heatid="70040" swimtime="00:00:30.48" reactiontime="+61" points="822">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="17" lane="7" heat="5" heatid="50004" swimtime="00:00:25.85" reactiontime="+57" points="838">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="304" place="17" lane="3" heat="1" heatid="10304" swimtime="00:00:25.78" reactiontime="+59" points="845">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="17" lane="1" heat="8" heatid="80030" swimtime="00:00:24.69" reactiontime="+60" points="801">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:24.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Turkmenistan" shortname="TKM" code="TKM" nation="TKM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="108075" lastname="ATAYEV" firstname="Merdan" gender="M" birthdate="1995-05-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.24" eventid="3" heat="2" lane="4">
                  <MEETINFO date="2021-07-25" />
                </ENTRY>
                <ENTRY entrytime="00:02:03.68" eventid="46" heat="1" lane="6">
                  <MEETINFO date="2021-07-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="34" lane="4" heat="2" heatid="20003" swimtime="00:00:55.04" reactiontime="+70" points="677">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.19" />
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                    <SPLIT distance="75" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:00:55.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="22" lane="6" heat="1" heatid="10046" swimtime="00:01:59.49" reactiontime="+70" points="690">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.76" />
                    <SPLIT distance="50" swimtime="00:00:28.23" />
                    <SPLIT distance="75" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:00:58.20" />
                    <SPLIT distance="125" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:28.75" />
                    <SPLIT distance="175" swimtime="00:01:44.30" />
                    <SPLIT distance="200" swimtime="00:01:59.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="118627" lastname="SEMYONOVA" firstname="Darya" gender="F" birthdate="2002-05-28">
              <ENTRIES>
                <ENTRY entrytime="00:01:01.31" eventid="13" heat="3" lane="4">
                  <MEETINFO date="2022-08-14" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="43" heat="1" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="50" lane="4" heat="3" heatid="30013" swimtime="00:00:59.20" reactiontime="+63" points="611">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.15" />
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                    <SPLIT distance="75" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:00:59.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="32" lane="1" heat="1" heatid="10043" swimtime="00:02:12.43" reactiontime="+64" points="577">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.93" />
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="75" swimtime="00:00:45.61" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="125" swimtime="00:01:19.72" />
                    <SPLIT distance="150" swimtime="00:01:37.40" />
                    <SPLIT distance="175" swimtime="00:01:55.03" />
                    <SPLIT distance="200" swimtime="00:02:12.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Timor-Leste" shortname="TLS" code="TLS" nation="TLS" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="183584" lastname="GUTERRES" firstname="Jolanio" gender="M" birthdate="2005-05-12">
              <ENTRIES>
                <ENTRY entrytime="00:01:11.08" eventid="14" heat="1" lane="6">
                  <MEETINFO date="2022-05-15" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.86" eventid="31" heat="2" lane="3">
                  <MEETINFO date="2022-05-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="84" lane="6" heat="1" heatid="10014" swimtime="00:01:10.23" reactiontime="+75" points="260">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.85" />
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                    <SPLIT distance="75" swimtime="00:00:50.34" />
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="76" lane="3" heat="2" heatid="20031" swimtime="00:00:29.09" reactiontime="+69" points="332">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110372" lastname="XIMENES BELO" firstname="Imelda" gender="F" birthdate="1998-10-24">
              <ENTRIES>
                <ENTRY entrytime="00:01:13.45" eventid="13" heat="2" lane="6">
                  <MEETINFO date="2022-05-14" />
                </ENTRY>
                <ENTRY entrytime="00:00:32.84" eventid="30" heat="2" lane="2">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="63" lane="6" heat="2" heatid="20013" swimtime="00:01:12.57" reactiontime="+76" points="331">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.62" />
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="75" swimtime="00:00:53.72" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="56" lane="2" heat="2" heatid="20030" swimtime="00:00:32.95" reactiontime="+54" points="337">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.03" />
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Togo" shortname="TOG" code="TOG" nation="TOG" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="209202" lastname="DAOU" firstname="Magnim Jordano" gender="M" birthdate="2004-07-11">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.60" eventid="5" heat="2" lane="5">
                  <MEETINFO date="2022-10-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:31.33" eventid="31" heat="2" lane="2">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="66" lane="5" heat="2" heatid="20005" swimtime="00:00:34.76" reactiontime="+70" points="244">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="78" lane="2" heat="2" heatid="20031" swimtime="00:00:30.39" reactiontime="+71" points="291">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.51" />
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197618" lastname="AMENOU" firstname="Marie" gender="F" birthdate="2006-08-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:43.73" eventid="4" heat="2" lane="8">
                  <MEETINFO date="2022-09-01" />
                </ENTRY>
                <ENTRY entrytime="00:00:34.58" eventid="30" heat="2" lane="7">
                  <MEETINFO date="2022-09-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="42" lane="8" heat="2" heatid="20004" swimtime="00:00:43.54" reactiontime="+78" points="175">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.87" />
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="57" lane="7" heat="2" heatid="20030" swimtime="00:00:34.70" reactiontime="+76" points="288">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Chinese Taipei" shortname="TPE" code="TPE" nation="TPE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="151877" lastname="CHUANG" firstname="Mu-Lun" gender="M" birthdate="2001-02-06">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.57" eventid="3" heat="2" lane="6">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="00:02:01.96" eventid="46" heat="1" lane="3">
                  <MEETINFO date="2022-03-10" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:25.55" eventid="19" heat="2" lane="7">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="29" lane="6" heat="2" heatid="20003" swimtime="00:00:52.79" reactiontime="+66" points="767">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.18" />
                    <SPLIT distance="50" swimtime="00:00:25.22" />
                    <SPLIT distance="75" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:00:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="-1" lane="3" heat="1" heatid="10046" swimtime="NT" status="DNS" />
                <RESULT eventid="19" place="27" lane="7" heat="2" heatid="20019" swimtime="00:00:24.15" reactiontime="+61" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                    <SPLIT distance="50" swimtime="00:00:24.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="101996" lastname="CAI" firstname="Bing Rong" gender="M" birthdate="1996-12-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.75" eventid="16" heat="2" lane="3">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="00:02:13.80" eventid="29" heat="2" lane="8">
                  <MEETINFO date="2021-09-17" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="40" lane="3" heat="2" heatid="20016" swimtime="00:01:00.16" reactiontime="+64" points="775">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.88" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:43.95" />
                    <SPLIT distance="100" swimtime="00:01:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="26" lane="8" heat="2" heatid="20029" swimtime="00:02:11.66" reactiontime="+64" points="760">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.34" />
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="75" swimtime="00:00:46.35" />
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                    <SPLIT distance="125" swimtime="00:01:20.38" />
                    <SPLIT distance="150" swimtime="00:01:37.47" />
                    <SPLIT distance="175" swimtime="00:01:54.63" />
                    <SPLIT distance="200" swimtime="00:02:11.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="154699" lastname="WANG" firstname="Kuan-Hung" gender="M" birthdate="2002-01-23">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.18" eventid="39" heat="5" lane="5">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="00:01:51.04" eventid="21" heat="2" lane="3">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="00:00:23.58" eventid="5" heat="5" lane="2">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="25" lane="5" heat="5" heatid="50039" swimtime="00:00:51.39" reactiontime="+56" points="803">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.13" />
                    <SPLIT distance="50" swimtime="00:00:23.80" />
                    <SPLIT distance="75" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="10" lane="3" heat="2" heatid="20021" swimtime="00:01:51.26" reactiontime="+57" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.53" />
                    <SPLIT distance="50" swimtime="00:00:25.52" />
                    <SPLIT distance="75" swimtime="00:00:39.63" />
                    <SPLIT distance="100" swimtime="00:00:54.11" />
                    <SPLIT distance="125" swimtime="00:01:08.76" />
                    <SPLIT distance="150" swimtime="00:01:22.98" />
                    <SPLIT distance="175" swimtime="00:01:37.18" />
                    <SPLIT distance="200" swimtime="00:01:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="47" lane="2" heat="5" heatid="50005" swimtime="00:00:23.68" reactiontime="+57" points="774">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.09" />
                    <SPLIT distance="50" swimtime="00:00:23.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156438" lastname="WANG" firstname="Hsing-Hao" gender="M" birthdate="1999-06-05">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.72" eventid="7" heat="2" lane="6">
                  <MEETINFO date="2021-07-28" />
                </ENTRY>
                <ENTRY entrytime="00:04:19.06" eventid="37" heat="1" lane="2">
                  <MEETINFO date="2021-07-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:54.19" eventid="23" heat="3" lane="8">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="7" place="26" lane="6" heat="2" heatid="20007" swimtime="00:01:58.57" reactiontime="+62" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.72" />
                    <SPLIT distance="50" swimtime="00:00:25.56" />
                    <SPLIT distance="75" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:00:56.31" />
                    <SPLIT distance="125" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:30.30" />
                    <SPLIT distance="175" swimtime="00:01:45.12" />
                    <SPLIT distance="200" swimtime="00:01:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="12" lane="2" heat="1" heatid="10037" swimtime="00:04:09.74" reactiontime="+60" points="831">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                    <SPLIT distance="75" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:00:57.73" />
                    <SPLIT distance="125" swimtime="00:01:14.31" />
                    <SPLIT distance="150" swimtime="00:01:30.03" />
                    <SPLIT distance="175" swimtime="00:01:46.23" />
                    <SPLIT distance="200" swimtime="00:02:02.32" />
                    <SPLIT distance="225" swimtime="00:02:19.84" />
                    <SPLIT distance="250" swimtime="00:02:37.39" />
                    <SPLIT distance="275" swimtime="00:02:54.96" />
                    <SPLIT distance="300" swimtime="00:03:12.79" />
                    <SPLIT distance="325" swimtime="00:03:27.67" />
                    <SPLIT distance="350" swimtime="00:03:41.90" />
                    <SPLIT distance="375" swimtime="00:03:56.05" />
                    <SPLIT distance="400" swimtime="00:04:09.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="-1" lane="8" heat="3" heatid="30023" swimtime="00:00:53.72" status="DSQ" reactiontime="+59" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="129429" lastname="WU" firstname="Chun-Feng" gender="M" birthdate="1990-12-02">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:28.34" eventid="41" heat="4" lane="7">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.88" eventid="31" heat="5" lane="3">
                  <MEETINFO date="2022-03-10" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="19" lane="7" heat="4" heatid="40041" swimtime="00:00:26.67" reactiontime="+67" points="818">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:26.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="45" lane="3" heat="5" heatid="50031" swimtime="00:00:22.05" reactiontime="+66" points="764">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.40" />
                    <SPLIT distance="50" swimtime="00:00:22.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156446" lastname="CHEN" firstname="Szu-An" gender="F" birthdate="2000-10-20">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:02:13.76" eventid="6" heat="2" lane="6">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="36" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="6" place="30" lane="6" heat="2" heatid="20006" swimtime="00:02:13.87" reactiontime="+72" points="754">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.27" />
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                    <SPLIT distance="75" swimtime="00:00:46.43" />
                    <SPLIT distance="100" swimtime="00:01:03.07" />
                    <SPLIT distance="125" swimtime="00:01:23.02" />
                    <SPLIT distance="150" swimtime="00:01:43.02" />
                    <SPLIT distance="175" swimtime="00:01:59.01" />
                    <SPLIT distance="200" swimtime="00:02:13.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="19" lane="3" heat="1" heatid="10036" swimtime="00:04:44.97" reactiontime="+69" points="750">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.91" />
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="75" swimtime="00:00:47.26" />
                    <SPLIT distance="100" swimtime="00:01:04.63" />
                    <SPLIT distance="125" swimtime="00:01:23.00" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                    <SPLIT distance="175" swimtime="00:01:59.58" />
                    <SPLIT distance="200" swimtime="00:02:18.72" />
                    <SPLIT distance="225" swimtime="00:02:37.95" />
                    <SPLIT distance="250" swimtime="00:02:58.50" />
                    <SPLIT distance="275" swimtime="00:03:19.07" />
                    <SPLIT distance="300" swimtime="00:03:39.81" />
                    <SPLIT distance="325" swimtime="00:03:56.34" />
                    <SPLIT distance="350" swimtime="00:04:12.53" />
                    <SPLIT distance="375" swimtime="00:04:29.14" />
                    <SPLIT distance="400" swimtime="00:04:44.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="157067" lastname="HUANG" firstname="Mei-Chien" gender="F" birthdate="1998-06-13">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:27.20" eventid="4" heat="3" lane="5">
                  <MEETINFO date="2022-06-23" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.99" eventid="30" heat="4" lane="3">
                  <MEETINFO date="2021-07-30" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="4" place="25" lane="5" heat="3" heatid="30004" swimtime="00:00:26.47" reactiontime="+65" points="781">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.16" />
                    <SPLIT distance="50" swimtime="00:00:26.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="25" lane="3" heat="4" heatid="40030" swimtime="00:00:25.07" reactiontime="+68" points="765">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:25.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213081" lastname="KUO" firstname="Jui-An" gender="F" birthdate="2005-02-01">
              <ENTRIES>
                <ENTRY entrytime="00:09:00.82" eventid="12" heat="1" lane="6">
                  <MEETINFO date="2022-07-15" />
                </ENTRY>
                <ENTRY entrytime="00:17:07.26" eventid="33" heat="1" lane="4">
                  <MEETINFO date="2022-07-15" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="19" lane="6" heat="1" heatid="10012" swimtime="00:09:01.45" reactiontime="+71" points="693">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="75" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:03.52" />
                    <SPLIT distance="125" swimtime="00:01:20.32" />
                    <SPLIT distance="150" swimtime="00:01:37.14" />
                    <SPLIT distance="175" swimtime="00:01:54.14" />
                    <SPLIT distance="200" swimtime="00:02:11.22" />
                    <SPLIT distance="225" swimtime="00:02:27.99" />
                    <SPLIT distance="250" swimtime="00:02:44.92" />
                    <SPLIT distance="275" swimtime="00:03:01.87" />
                    <SPLIT distance="300" swimtime="00:03:19.09" />
                    <SPLIT distance="325" swimtime="00:03:36.23" />
                    <SPLIT distance="350" swimtime="00:03:53.64" />
                    <SPLIT distance="375" swimtime="00:04:10.72" />
                    <SPLIT distance="400" swimtime="00:04:27.95" />
                    <SPLIT distance="425" swimtime="00:04:45.00" />
                    <SPLIT distance="450" swimtime="00:05:02.19" />
                    <SPLIT distance="475" swimtime="00:05:19.18" />
                    <SPLIT distance="500" swimtime="00:05:36.24" />
                    <SPLIT distance="525" swimtime="00:05:53.17" />
                    <SPLIT distance="550" swimtime="00:06:10.21" />
                    <SPLIT distance="575" swimtime="00:06:27.38" />
                    <SPLIT distance="600" swimtime="00:06:44.56" />
                    <SPLIT distance="625" swimtime="00:07:01.75" />
                    <SPLIT distance="650" swimtime="00:07:19.07" />
                    <SPLIT distance="675" swimtime="00:07:36.14" />
                    <SPLIT distance="700" swimtime="00:07:53.46" />
                    <SPLIT distance="725" swimtime="00:08:10.62" />
                    <SPLIT distance="750" swimtime="00:08:28.09" />
                    <SPLIT distance="775" swimtime="00:08:44.94" />
                    <SPLIT distance="800" swimtime="00:09:01.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="16" lane="4" heat="1" heatid="10033" swimtime="00:17:16.69" reactiontime="+50" points="694">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.76" />
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                    <SPLIT distance="75" swimtime="00:00:48.06" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="125" swimtime="00:01:21.77" />
                    <SPLIT distance="150" swimtime="00:01:38.85" />
                    <SPLIT distance="175" swimtime="00:01:55.85" />
                    <SPLIT distance="200" swimtime="00:02:12.85" />
                    <SPLIT distance="225" swimtime="00:02:29.90" />
                    <SPLIT distance="250" swimtime="00:02:47.06" />
                    <SPLIT distance="275" swimtime="00:03:04.09" />
                    <SPLIT distance="300" swimtime="00:03:21.25" />
                    <SPLIT distance="325" swimtime="00:03:38.27" />
                    <SPLIT distance="350" swimtime="00:03:55.54" />
                    <SPLIT distance="375" swimtime="00:04:12.59" />
                    <SPLIT distance="400" swimtime="00:04:29.78" />
                    <SPLIT distance="425" swimtime="00:04:47.06" />
                    <SPLIT distance="450" swimtime="00:05:04.14" />
                    <SPLIT distance="475" swimtime="00:05:21.37" />
                    <SPLIT distance="500" swimtime="00:05:38.70" />
                    <SPLIT distance="525" swimtime="00:05:55.87" />
                    <SPLIT distance="550" swimtime="00:06:13.26" />
                    <SPLIT distance="575" swimtime="00:06:30.53" />
                    <SPLIT distance="600" swimtime="00:06:48.17" />
                    <SPLIT distance="625" swimtime="00:07:05.60" />
                    <SPLIT distance="650" swimtime="00:07:23.09" />
                    <SPLIT distance="675" swimtime="00:07:40.60" />
                    <SPLIT distance="700" swimtime="00:07:58.22" />
                    <SPLIT distance="725" swimtime="00:08:15.80" />
                    <SPLIT distance="750" swimtime="00:08:33.49" />
                    <SPLIT distance="775" swimtime="00:08:51.04" />
                    <SPLIT distance="800" swimtime="00:09:08.57" />
                    <SPLIT distance="825" swimtime="00:09:26.15" />
                    <SPLIT distance="850" swimtime="00:09:43.64" />
                    <SPLIT distance="875" swimtime="00:10:01.15" />
                    <SPLIT distance="900" swimtime="00:10:18.63" />
                    <SPLIT distance="925" swimtime="00:10:35.87" />
                    <SPLIT distance="950" swimtime="00:10:53.48" />
                    <SPLIT distance="975" swimtime="00:11:10.85" />
                    <SPLIT distance="1000" swimtime="00:11:28.35" />
                    <SPLIT distance="1025" swimtime="00:11:45.72" />
                    <SPLIT distance="1050" swimtime="00:12:03.02" />
                    <SPLIT distance="1075" swimtime="00:12:20.19" />
                    <SPLIT distance="1100" swimtime="00:12:37.77" />
                    <SPLIT distance="1125" swimtime="00:12:55.24" />
                    <SPLIT distance="1150" swimtime="00:13:12.89" />
                    <SPLIT distance="1175" swimtime="00:13:30.53" />
                    <SPLIT distance="1200" swimtime="00:13:48.31" />
                    <SPLIT distance="1225" swimtime="00:14:06.13" />
                    <SPLIT distance="1250" swimtime="00:14:23.83" />
                    <SPLIT distance="1275" swimtime="00:14:41.33" />
                    <SPLIT distance="1300" swimtime="00:14:58.78" />
                    <SPLIT distance="1325" swimtime="00:15:16.14" />
                    <SPLIT distance="1350" swimtime="00:15:33.78" />
                    <SPLIT distance="1375" swimtime="00:15:51.30" />
                    <SPLIT distance="1400" swimtime="00:16:08.85" />
                    <SPLIT distance="1425" swimtime="00:16:26.19" />
                    <SPLIT distance="1450" swimtime="00:16:43.35" />
                    <SPLIT distance="1475" swimtime="00:17:00.37" />
                    <SPLIT distance="1500" swimtime="00:17:16.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Chinese Taipei">
              <RESULTS>
                <RESULT eventid="9" place="12" lane="1" heat="1" swimtime="00:03:17.25" reactiontime="+56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.79" />
                    <SPLIT distance="50" swimtime="00:00:22.79" />
                    <SPLIT distance="75" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:00:48.33" />
                    <SPLIT distance="125" swimtime="00:00:59.03" />
                    <SPLIT distance="150" swimtime="00:01:11.23" />
                    <SPLIT distance="175" swimtime="00:01:24.16" />
                    <SPLIT distance="200" swimtime="00:01:37.22" />
                    <SPLIT distance="225" swimtime="00:01:48.57" />
                    <SPLIT distance="250" swimtime="00:02:01.64" />
                    <SPLIT distance="275" swimtime="00:02:15.00" />
                    <SPLIT distance="300" swimtime="00:02:28.19" />
                    <SPLIT distance="325" swimtime="00:02:39.38" />
                    <SPLIT distance="350" swimtime="00:02:52.03" />
                    <SPLIT distance="375" swimtime="00:03:04.70" />
                    <SPLIT distance="400" swimtime="00:03:17.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154699" reactiontime="+56" />
                    <RELAYPOSITION number="2" athleteid="151877" reactiontime="+43" />
                    <RELAYPOSITION number="3" athleteid="101996" reactiontime="+45" />
                    <RELAYPOSITION number="4" athleteid="156438" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Chinese Taipei">
              <RESULTS>
                <RESULT eventid="48" place="-1" lane="4" heat="1" status="DNS" swimtime="NT" />
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Chinese Taipei">
              <RESULTS>
                <RESULT eventid="26" place="13" lane="6" heat="1" swimtime="00:01:30.09" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.43" />
                    <SPLIT distance="50" swimtime="00:00:22.22" />
                    <SPLIT distance="75" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:00:45.37" />
                    <SPLIT distance="125" swimtime="00:00:56.28" />
                    <SPLIT distance="150" swimtime="00:01:08.20" />
                    <SPLIT distance="175" swimtime="00:01:18.55" />
                    <SPLIT distance="200" swimtime="00:01:30.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="129429" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="101996" reactiontime="+31" />
                    <RELAYPOSITION number="3" athleteid="156438" reactiontime="+41" />
                    <RELAYPOSITION number="4" athleteid="151877" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Chinese Taipei">
              <RESULTS>
                <RESULT eventid="27" place="12" lane="8" heat="4" swimtime="00:01:34.87" reactiontime="+57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.87" />
                    <SPLIT distance="50" swimtime="00:00:22.47" />
                    <SPLIT distance="75" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:00:44.24" />
                    <SPLIT distance="125" swimtime="00:00:56.68" />
                    <SPLIT distance="150" swimtime="00:01:10.01" />
                    <SPLIT distance="175" swimtime="00:01:21.73" />
                    <SPLIT distance="200" swimtime="00:01:34.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="154699" reactiontime="+57" />
                    <RELAYPOSITION number="2" athleteid="129429" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="156446" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="157067" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Chinese Taipei">
              <RESULTS>
                <RESULT eventid="11" place="18" lane="6" heat="1" swimtime="00:01:43.48" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.04" />
                    <SPLIT distance="50" swimtime="00:00:24.57" />
                    <SPLIT distance="75" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:00:51.37" />
                    <SPLIT distance="125" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:17.58" />
                    <SPLIT distance="175" swimtime="00:01:30.00" />
                    <SPLIT distance="200" swimtime="00:01:43.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="151877" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="129429" reactiontime="+21" />
                    <RELAYPOSITION number="3" athleteid="157067" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="156446" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Chinese Taipei">
              <RESULTS>
                <RESULT eventid="35" place="-1" lane="6" heat="3" status="DSQ" swimtime="00:01:37.05" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:24.20" />
                    <SPLIT distance="75" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:00:50.57" />
                    <SPLIT distance="125" swimtime="00:01:01.24" />
                    <SPLIT distance="150" swimtime="00:01:13.97" />
                    <SPLIT distance="175" swimtime="00:01:25.05" />
                    <SPLIT distance="200" swimtime="00:01:37.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="151877" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="129429" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="154699" reactiontime="+24" status="DSQ" />
                    <RELAYPOSITION number="4" athleteid="156438" reactiontime="+40" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Trinidad &amp; Tobago" shortname="TTO" code="TTO" nation="TTO" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="118453" lastname="CARTER" firstname="Dylan" gender="M" birthdate="1996-01-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:22.72" eventid="19" heat="5" lane="4">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.98" eventid="5" heat="8" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:20.72" eventid="31" heat="9" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="119" place="7" lane="2" heat="1" heatid="10119" swimtime="00:00:23.12" reactiontime="+56" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="4" lane="4" heat="5" heatid="50019" swimtime="00:00:23.07" reactiontime="+52" points="893">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:23.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="5" lane="5" heat="1" heatid="10219" swimtime="00:00:22.90" reactiontime="+54" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:22.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="105" place="6" lane="5" heat="1" heatid="10105" swimtime="00:00:22.14" reactiontime="+62" points="948">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.10" />
                    <SPLIT distance="50" swimtime="00:00:22.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="4" lane="4" heat="8" heatid="80005" swimtime="00:00:22.11" reactiontime="+61" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.01" />
                    <SPLIT distance="50" swimtime="00:00:22.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="2" lane="5" heat="1" heatid="10205" swimtime="00:00:22.02" reactiontime="+62" points="963">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.02" />
                    <SPLIT distance="50" swimtime="00:00:22.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="131" place="3" lane="7" heat="1" heatid="10131" swimtime="00:00:20.72" reactiontime="+61" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.05" />
                    <SPLIT distance="50" swimtime="00:00:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="2" lane="4" heat="9" heatid="90031" swimtime="00:00:20.70" reactiontime="+63" points="923">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.03" />
                    <SPLIT distance="50" swimtime="00:00:20.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="5" lane="4" heat="1" heatid="10231" swimtime="00:00:20.94" reactiontime="+62" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.06" />
                    <SPLIT distance="50" swimtime="00:00:20.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Tunisia" shortname="TUN" code="TUN" nation="TUN" type="NOC">
          <ATHLETES />
        </CLUB>
        <CLUB name="Turkey" shortname="TUR" code="TUR" nation="TUR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197192" lastname="GOR" firstname="Rasim Ogulcan" gender="M" birthdate="1998-10-19">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.92" eventid="3" heat="6" lane="8">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.62" eventid="19" heat="6" lane="1">
                  <MEETINFO date="2021-12-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="27" lane="8" heat="6" heatid="60003" swimtime="00:00:52.54" reactiontime="+63" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="75" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="28" lane="1" heat="6" heatid="60019" swimtime="00:00:24.29" reactiontime="+62" points="765">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:24.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110514" lastname="SAKCI" firstname="Huseyin" gender="M" birthdate="1997-11-15">
              <ENTRIES>
                <ENTRY entrytime="00:00:56.25" eventid="16" heat="8" lane="5">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.38" eventid="41" heat="8" lane="4">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.36" eventid="31" heat="10" lane="1">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:00:54.60" eventid="23" heat="2" lane="6">
                  <MEETINFO date="2022-10-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="13" lane="5" heat="8" heatid="80016" swimtime="00:00:57.70" reactiontime="+66" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="75" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:00:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="12" lane="1" heat="2" heatid="20216" swimtime="00:00:57.65" reactiontime="+64" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                    <SPLIT distance="75" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:00:57.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="8" lane="8" heat="1" heatid="10141" swimtime="00:00:26.09" reactiontime="+64" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.73" />
                    <SPLIT distance="50" swimtime="00:00:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="9" lane="4" heat="8" heatid="80041" swimtime="00:00:26.26" reactiontime="+68" points="857">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:26.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="8" lane="2" heat="2" heatid="20241" swimtime="00:00:26.04" reactiontime="+64" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="39" lane="1" heat="10" heatid="100031" swimtime="00:00:21.65" reactiontime="+64" points="807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.41" />
                    <SPLIT distance="50" swimtime="00:00:21.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="17" lane="6" heat="2" heatid="20023" swimtime="00:00:52.81" reactiontime="+68" points="812">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.57" />
                    <SPLIT distance="50" swimtime="00:00:24.48" />
                    <SPLIT distance="75" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:00:52.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="323" place="17" lane="4" heat="1" heatid="10323" swimtime="00:00:52.24" reactiontime="+62" points="839">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:24.44" />
                    <SPLIT distance="75" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:00:52.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156135" lastname="OGRETIR" firstname="Berkay" gender="M" birthdate="1998-02-16">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.17" eventid="16" heat="6" lane="6">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:02:06.75" eventid="29" heat="5" lane="1">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="26" lane="6" heat="6" heatid="60016" swimtime="00:00:58.27" reactiontime="+64" points="853">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.62" />
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                    <SPLIT distance="75" swimtime="00:00:42.61" />
                    <SPLIT distance="100" swimtime="00:00:58.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="17" lane="1" heat="5" heatid="50029" swimtime="00:02:07.12" reactiontime="+68" points="844">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                    <SPLIT distance="75" swimtime="00:00:44.28" />
                    <SPLIT distance="100" swimtime="00:01:00.13" />
                    <SPLIT distance="125" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:32.83" />
                    <SPLIT distance="175" swimtime="00:01:49.67" />
                    <SPLIT distance="200" swimtime="00:02:07.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150083" lastname="GURES" firstname="Umitcan" gender="M" birthdate="1999-06-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.80" eventid="39" heat="6" lane="6">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.37" eventid="5" heat="9" lane="6">
                  <MEETINFO date="2021-11-06" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="35" lane="6" heat="6" heatid="60039" swimtime="00:00:52.94" reactiontime="+60" points="735">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.14" />
                    <SPLIT distance="50" swimtime="00:00:24.46" />
                    <SPLIT distance="75" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:00:52.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="21" lane="6" heat="9" heatid="90005" swimtime="00:00:22.75" reactiontime="+60" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.55" />
                    <SPLIT distance="50" swimtime="00:00:22.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170692" lastname="KILAVUZ" firstname="Mert" gender="M" birthdate="2003-08-26">
              <ENTRIES>
                <ENTRY entrytime="00:03:55.70" eventid="24" heat="1" lane="4">
                  <MEETINFO date="2022-05-15" />
                </ENTRY>
                <ENTRY entrytime="00:07:43.64" eventid="42" heat="2" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="24" place="21" lane="4" heat="1" heatid="10024" swimtime="00:03:46.32" reactiontime="+76" points="824">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.50" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                    <SPLIT distance="75" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:00:54.11" />
                    <SPLIT distance="125" swimtime="00:01:08.14" />
                    <SPLIT distance="150" swimtime="00:01:22.43" />
                    <SPLIT distance="175" swimtime="00:01:36.70" />
                    <SPLIT distance="200" swimtime="00:01:51.19" />
                    <SPLIT distance="225" swimtime="00:02:05.58" />
                    <SPLIT distance="250" swimtime="00:02:20.00" />
                    <SPLIT distance="275" swimtime="00:02:34.47" />
                    <SPLIT distance="300" swimtime="00:02:48.99" />
                    <SPLIT distance="325" swimtime="00:03:03.45" />
                    <SPLIT distance="350" swimtime="00:03:18.13" />
                    <SPLIT distance="375" swimtime="00:03:32.43" />
                    <SPLIT distance="400" swimtime="00:03:46.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="13" lane="4" heat="2" heatid="20042" swimtime="00:07:47.57" reactiontime="+74" points="852">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.85" />
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                    <SPLIT distance="75" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:00:55.95" />
                    <SPLIT distance="125" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:25.10" />
                    <SPLIT distance="175" swimtime="00:01:39.71" />
                    <SPLIT distance="200" swimtime="00:01:54.35" />
                    <SPLIT distance="225" swimtime="00:02:08.96" />
                    <SPLIT distance="250" swimtime="00:02:23.60" />
                    <SPLIT distance="275" swimtime="00:02:38.16" />
                    <SPLIT distance="300" swimtime="00:02:52.80" />
                    <SPLIT distance="325" swimtime="00:03:07.43" />
                    <SPLIT distance="350" swimtime="00:03:22.22" />
                    <SPLIT distance="375" swimtime="00:03:36.95" />
                    <SPLIT distance="400" swimtime="00:03:51.83" />
                    <SPLIT distance="425" swimtime="00:04:06.63" />
                    <SPLIT distance="450" swimtime="00:04:21.45" />
                    <SPLIT distance="475" swimtime="00:04:36.22" />
                    <SPLIT distance="500" swimtime="00:04:51.19" />
                    <SPLIT distance="525" swimtime="00:05:05.97" />
                    <SPLIT distance="550" swimtime="00:05:20.84" />
                    <SPLIT distance="575" swimtime="00:05:35.60" />
                    <SPLIT distance="600" swimtime="00:05:50.51" />
                    <SPLIT distance="625" swimtime="00:06:05.41" />
                    <SPLIT distance="650" swimtime="00:06:20.28" />
                    <SPLIT distance="675" swimtime="00:06:35.03" />
                    <SPLIT distance="700" swimtime="00:06:49.80" />
                    <SPLIT distance="725" swimtime="00:07:04.45" />
                    <SPLIT distance="750" swimtime="00:07:19.27" />
                    <SPLIT distance="775" swimtime="00:07:33.72" />
                    <SPLIT distance="800" swimtime="00:07:47.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="122443" lastname="TEKIN" firstname="Doruk" gender="M" birthdate="1994-12-21">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:23.54" eventid="19" heat="6" lane="7">
                  <MEETINFO date="2021-11-02" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="19" place="32" lane="7" heat="6" heatid="60019" swimtime="00:00:24.63" reactiontime="+59" points="734">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.96" />
                    <SPLIT distance="50" swimtime="00:00:24.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="110602" lastname="USTUNDAG" firstname="Nida" gender="F" birthdate="1996-10-21">
              <ENTRIES>
                <ENTRY entrytime="00:02:08.14" eventid="20" heat="4" lane="7">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="20" place="15" lane="7" heat="4" heatid="40020" swimtime="00:02:09.14" reactiontime="+74" points="794">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                    <SPLIT distance="75" swimtime="00:00:45.43" />
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                    <SPLIT distance="125" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:01:34.78" />
                    <SPLIT distance="175" swimtime="00:01:51.61" />
                    <SPLIT distance="200" swimtime="00:02:09.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170682" lastname="TUNCEL" firstname="Merve" gender="F" birthdate="2005-01-01">
              <ENTRIES>
                <ENTRY entrytime="00:02:00.02" eventid="43" heat="2" lane="3">
                  <MEETINFO date="2022-07-06" />
                </ENTRY>
                <ENTRY entrytime="00:04:02.47" eventid="1" heat="3" lane="2">
                  <MEETINFO date="2021-11-07" />
                </ENTRY>
                <ENTRY entrytime="00:08:17.12" eventid="12" heat="0" lane="2147483647">
                  <MEETINFO date="2021-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="00:15:50.36" eventid="33" heat="0" lane="2147483647">
                  <MEETINFO date="2021-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="23" lane="3" heat="2" heatid="20043" swimtime="00:01:59.32" reactiontime="+68" points="790">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="75" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:00:58.45" />
                    <SPLIT distance="125" swimtime="00:01:13.62" />
                    <SPLIT distance="150" swimtime="00:01:28.98" />
                    <SPLIT distance="175" swimtime="00:01:44.32" />
                    <SPLIT distance="200" swimtime="00:01:59.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="17" lane="2" heat="3" heatid="30001" swimtime="00:04:10.60" reactiontime="+69" points="813">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.89" />
                    <SPLIT distance="50" swimtime="00:00:29.03" />
                    <SPLIT distance="75" swimtime="00:00:44.40" />
                    <SPLIT distance="100" swimtime="00:00:59.89" />
                    <SPLIT distance="125" swimtime="00:01:15.39" />
                    <SPLIT distance="150" swimtime="00:01:31.04" />
                    <SPLIT distance="175" swimtime="00:01:46.63" />
                    <SPLIT distance="200" swimtime="00:02:02.51" />
                    <SPLIT distance="225" swimtime="00:02:18.36" />
                    <SPLIT distance="250" swimtime="00:02:34.33" />
                    <SPLIT distance="275" swimtime="00:02:50.36" />
                    <SPLIT distance="300" swimtime="00:03:06.48" />
                    <SPLIT distance="325" swimtime="00:03:22.59" />
                    <SPLIT distance="350" swimtime="00:03:38.77" />
                    <SPLIT distance="375" swimtime="00:03:54.89" />
                    <SPLIT distance="400" swimtime="00:04:10.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="5" lane="2" heat="5" heatid="30112" swimtime="00:08:17.89" reactiontime="+68" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                    <SPLIT distance="75" swimtime="00:00:44.19" />
                    <SPLIT distance="100" swimtime="00:00:59.68" />
                    <SPLIT distance="125" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:30.78" />
                    <SPLIT distance="175" swimtime="00:01:46.32" />
                    <SPLIT distance="200" swimtime="00:02:01.89" />
                    <SPLIT distance="225" swimtime="00:02:17.44" />
                    <SPLIT distance="250" swimtime="00:02:33.07" />
                    <SPLIT distance="275" swimtime="00:02:48.60" />
                    <SPLIT distance="300" swimtime="00:03:04.37" />
                    <SPLIT distance="325" swimtime="00:03:19.96" />
                    <SPLIT distance="350" swimtime="00:03:35.77" />
                    <SPLIT distance="375" swimtime="00:03:51.40" />
                    <SPLIT distance="400" swimtime="00:04:07.22" />
                    <SPLIT distance="425" swimtime="00:04:22.90" />
                    <SPLIT distance="450" swimtime="00:04:38.59" />
                    <SPLIT distance="475" swimtime="00:04:54.34" />
                    <SPLIT distance="500" swimtime="00:05:10.02" />
                    <SPLIT distance="525" swimtime="00:05:25.78" />
                    <SPLIT distance="550" swimtime="00:05:41.46" />
                    <SPLIT distance="575" swimtime="00:05:57.25" />
                    <SPLIT distance="600" swimtime="00:06:12.88" />
                    <SPLIT distance="625" swimtime="00:06:28.48" />
                    <SPLIT distance="650" swimtime="00:06:44.12" />
                    <SPLIT distance="675" swimtime="00:06:59.86" />
                    <SPLIT distance="700" swimtime="00:07:15.75" />
                    <SPLIT distance="725" swimtime="00:07:31.56" />
                    <SPLIT distance="750" swimtime="00:07:47.26" />
                    <SPLIT distance="775" swimtime="00:08:03.05" />
                    <SPLIT distance="800" swimtime="00:08:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="7" lane="5" heat="5" heatid="30133" swimtime="00:15:58.05" reactiontime="+69" points="879">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.05" />
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                    <SPLIT distance="75" swimtime="00:00:44.58" />
                    <SPLIT distance="100" swimtime="00:01:00.18" />
                    <SPLIT distance="125" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:31.58" />
                    <SPLIT distance="175" swimtime="00:01:47.31" />
                    <SPLIT distance="200" swimtime="00:02:02.99" />
                    <SPLIT distance="225" swimtime="00:02:18.66" />
                    <SPLIT distance="250" swimtime="00:02:34.40" />
                    <SPLIT distance="275" swimtime="00:02:50.32" />
                    <SPLIT distance="300" swimtime="00:03:06.13" />
                    <SPLIT distance="325" swimtime="00:03:21.86" />
                    <SPLIT distance="350" swimtime="00:03:37.68" />
                    <SPLIT distance="375" swimtime="00:03:53.62" />
                    <SPLIT distance="400" swimtime="00:04:09.44" />
                    <SPLIT distance="425" swimtime="00:04:25.21" />
                    <SPLIT distance="450" swimtime="00:04:41.09" />
                    <SPLIT distance="475" swimtime="00:04:57.02" />
                    <SPLIT distance="500" swimtime="00:05:12.88" />
                    <SPLIT distance="525" swimtime="00:05:28.82" />
                    <SPLIT distance="550" swimtime="00:05:44.78" />
                    <SPLIT distance="575" swimtime="00:06:00.79" />
                    <SPLIT distance="600" swimtime="00:06:16.71" />
                    <SPLIT distance="625" swimtime="00:06:32.74" />
                    <SPLIT distance="650" swimtime="00:06:48.64" />
                    <SPLIT distance="675" swimtime="00:07:04.60" />
                    <SPLIT distance="700" swimtime="00:07:20.65" />
                    <SPLIT distance="725" swimtime="00:07:36.61" />
                    <SPLIT distance="750" swimtime="00:07:52.66" />
                    <SPLIT distance="775" swimtime="00:08:08.73" />
                    <SPLIT distance="800" swimtime="00:08:24.78" />
                    <SPLIT distance="825" swimtime="00:08:40.83" />
                    <SPLIT distance="850" swimtime="00:08:56.99" />
                    <SPLIT distance="875" swimtime="00:09:13.02" />
                    <SPLIT distance="900" swimtime="00:09:29.11" />
                    <SPLIT distance="925" swimtime="00:09:45.28" />
                    <SPLIT distance="950" swimtime="00:10:01.39" />
                    <SPLIT distance="975" swimtime="00:10:17.54" />
                    <SPLIT distance="1000" swimtime="00:10:33.47" />
                    <SPLIT distance="1025" swimtime="00:10:49.70" />
                    <SPLIT distance="1050" swimtime="00:11:05.84" />
                    <SPLIT distance="1075" swimtime="00:11:22.05" />
                    <SPLIT distance="1100" swimtime="00:11:38.20" />
                    <SPLIT distance="1125" swimtime="00:11:54.39" />
                    <SPLIT distance="1150" swimtime="00:12:10.65" />
                    <SPLIT distance="1175" swimtime="00:12:26.73" />
                    <SPLIT distance="1200" swimtime="00:12:42.87" />
                    <SPLIT distance="1225" swimtime="00:12:59.04" />
                    <SPLIT distance="1250" swimtime="00:13:15.18" />
                    <SPLIT distance="1275" swimtime="00:13:31.29" />
                    <SPLIT distance="1300" swimtime="00:13:47.39" />
                    <SPLIT distance="1325" swimtime="00:14:03.49" />
                    <SPLIT distance="1350" swimtime="00:14:19.42" />
                    <SPLIT distance="1375" swimtime="00:14:35.52" />
                    <SPLIT distance="1400" swimtime="00:14:51.82" />
                    <SPLIT distance="1425" swimtime="00:15:08.31" />
                    <SPLIT distance="1450" swimtime="00:15:24.99" />
                    <SPLIT distance="1475" swimtime="00:15:41.69" />
                    <SPLIT distance="1500" swimtime="00:15:58.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="170684" lastname="ERTAN" firstname="Deniz" gender="F" birthdate="2004-01-01">
              <ENTRIES>
                <ENTRY entrytime="00:04:40.45" eventid="36" heat="2" lane="3">
                  <MEETINFO date="2022-04-13" />
                </ENTRY>
                <ENTRY entrytime="00:08:24.94" eventid="12" heat="2" lane="5">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="00:15:51.65" eventid="33" heat="0" lane="2147483647">
                  <MEETINFO date="2021-11-04" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="36" place="13" lane="3" heat="2" heatid="20036" swimtime="00:04:38.11" reactiontime="+70" points="807">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="75" swimtime="00:00:46.31" />
                    <SPLIT distance="100" swimtime="00:01:03.23" />
                    <SPLIT distance="125" swimtime="00:01:22.16" />
                    <SPLIT distance="150" swimtime="00:01:40.35" />
                    <SPLIT distance="175" swimtime="00:01:58.49" />
                    <SPLIT distance="200" swimtime="00:02:16.62" />
                    <SPLIT distance="225" swimtime="00:02:35.75" />
                    <SPLIT distance="250" swimtime="00:02:55.07" />
                    <SPLIT distance="275" swimtime="00:03:14.71" />
                    <SPLIT distance="300" swimtime="00:03:34.41" />
                    <SPLIT distance="325" swimtime="00:03:51.16" />
                    <SPLIT distance="350" swimtime="00:04:07.06" />
                    <SPLIT distance="375" swimtime="00:04:22.86" />
                    <SPLIT distance="400" swimtime="00:04:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="11" lane="5" heat="2" heatid="20012" swimtime="00:08:29.92" reactiontime="+70" points="830">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.67" />
                    <SPLIT distance="50" swimtime="00:00:28.74" />
                    <SPLIT distance="75" swimtime="00:00:44.13" />
                    <SPLIT distance="100" swimtime="00:00:59.96" />
                    <SPLIT distance="125" swimtime="00:01:15.60" />
                    <SPLIT distance="150" swimtime="00:01:31.43" />
                    <SPLIT distance="175" swimtime="00:01:47.25" />
                    <SPLIT distance="200" swimtime="00:02:03.35" />
                    <SPLIT distance="225" swimtime="00:02:19.13" />
                    <SPLIT distance="250" swimtime="00:02:35.18" />
                    <SPLIT distance="275" swimtime="00:02:51.08" />
                    <SPLIT distance="300" swimtime="00:03:07.12" />
                    <SPLIT distance="325" swimtime="00:03:23.08" />
                    <SPLIT distance="350" swimtime="00:03:39.24" />
                    <SPLIT distance="375" swimtime="00:03:55.14" />
                    <SPLIT distance="400" swimtime="00:04:11.28" />
                    <SPLIT distance="425" swimtime="00:04:27.29" />
                    <SPLIT distance="450" swimtime="00:04:43.49" />
                    <SPLIT distance="475" swimtime="00:04:59.50" />
                    <SPLIT distance="500" swimtime="00:05:15.71" />
                    <SPLIT distance="525" swimtime="00:05:31.71" />
                    <SPLIT distance="550" swimtime="00:05:47.96" />
                    <SPLIT distance="575" swimtime="00:06:04.13" />
                    <SPLIT distance="600" swimtime="00:06:20.45" />
                    <SPLIT distance="625" swimtime="00:06:36.65" />
                    <SPLIT distance="650" swimtime="00:06:53.14" />
                    <SPLIT distance="675" swimtime="00:07:09.40" />
                    <SPLIT distance="700" swimtime="00:07:25.76" />
                    <SPLIT distance="725" swimtime="00:07:41.89" />
                    <SPLIT distance="750" swimtime="00:07:58.25" />
                    <SPLIT distance="775" swimtime="00:08:14.30" />
                    <SPLIT distance="800" swimtime="00:08:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="6" lane="3" heat="5" heatid="30133" swimtime="00:15:53.73" reactiontime="+71" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="75" swimtime="00:00:44.50" />
                    <SPLIT distance="100" swimtime="00:01:00.24" />
                    <SPLIT distance="125" swimtime="00:01:15.92" />
                    <SPLIT distance="150" swimtime="00:01:31.68" />
                    <SPLIT distance="175" swimtime="00:01:47.47" />
                    <SPLIT distance="200" swimtime="00:02:03.41" />
                    <SPLIT distance="225" swimtime="00:02:19.22" />
                    <SPLIT distance="250" swimtime="00:02:35.06" />
                    <SPLIT distance="275" swimtime="00:02:51.04" />
                    <SPLIT distance="300" swimtime="00:03:06.83" />
                    <SPLIT distance="325" swimtime="00:03:22.68" />
                    <SPLIT distance="350" swimtime="00:03:38.53" />
                    <SPLIT distance="375" swimtime="00:03:54.40" />
                    <SPLIT distance="400" swimtime="00:04:10.24" />
                    <SPLIT distance="425" swimtime="00:04:26.11" />
                    <SPLIT distance="450" swimtime="00:04:42.08" />
                    <SPLIT distance="475" swimtime="00:04:58.01" />
                    <SPLIT distance="500" swimtime="00:05:13.96" />
                    <SPLIT distance="525" swimtime="00:05:29.98" />
                    <SPLIT distance="550" swimtime="00:05:45.91" />
                    <SPLIT distance="575" swimtime="00:06:01.88" />
                    <SPLIT distance="600" swimtime="00:06:17.88" />
                    <SPLIT distance="625" swimtime="00:06:33.82" />
                    <SPLIT distance="650" swimtime="00:06:49.90" />
                    <SPLIT distance="675" swimtime="00:07:05.97" />
                    <SPLIT distance="700" swimtime="00:07:22.00" />
                    <SPLIT distance="725" swimtime="00:07:38.04" />
                    <SPLIT distance="750" swimtime="00:07:54.16" />
                    <SPLIT distance="775" swimtime="00:08:10.18" />
                    <SPLIT distance="800" swimtime="00:08:26.17" />
                    <SPLIT distance="825" swimtime="00:08:42.22" />
                    <SPLIT distance="850" swimtime="00:08:58.35" />
                    <SPLIT distance="875" swimtime="00:09:14.46" />
                    <SPLIT distance="900" swimtime="00:09:30.44" />
                    <SPLIT distance="925" swimtime="00:09:46.37" />
                    <SPLIT distance="950" swimtime="00:10:02.45" />
                    <SPLIT distance="975" swimtime="00:10:18.65" />
                    <SPLIT distance="1000" swimtime="00:10:34.75" />
                    <SPLIT distance="1025" swimtime="00:10:50.78" />
                    <SPLIT distance="1050" swimtime="00:11:06.88" />
                    <SPLIT distance="1075" swimtime="00:11:23.04" />
                    <SPLIT distance="1100" swimtime="00:11:39.12" />
                    <SPLIT distance="1125" swimtime="00:11:55.12" />
                    <SPLIT distance="1150" swimtime="00:12:11.20" />
                    <SPLIT distance="1175" swimtime="00:12:27.11" />
                    <SPLIT distance="1200" swimtime="00:12:42.97" />
                    <SPLIT distance="1225" swimtime="00:12:58.90" />
                    <SPLIT distance="1250" swimtime="00:13:14.83" />
                    <SPLIT distance="1275" swimtime="00:13:30.86" />
                    <SPLIT distance="1300" swimtime="00:13:46.83" />
                    <SPLIT distance="1325" swimtime="00:14:02.80" />
                    <SPLIT distance="1350" swimtime="00:14:18.84" />
                    <SPLIT distance="1375" swimtime="00:14:34.88" />
                    <SPLIT distance="1400" swimtime="00:14:50.82" />
                    <SPLIT distance="1425" swimtime="00:15:06.72" />
                    <SPLIT distance="1450" swimtime="00:15:22.57" />
                    <SPLIT distance="1475" swimtime="00:15:38.46" />
                    <SPLIT distance="1500" swimtime="00:15:53.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Turkey">
              <RESULTS>
                <RESULT eventid="48" place="15" lane="2" heat="3" swimtime="00:03:34.89" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.33" />
                    <SPLIT distance="50" swimtime="00:00:25.94" />
                    <SPLIT distance="75" swimtime="00:00:40.38" />
                    <SPLIT distance="100" swimtime="00:00:55.10" />
                    <SPLIT distance="125" swimtime="00:01:07.12" />
                    <SPLIT distance="150" swimtime="00:01:21.85" />
                    <SPLIT distance="175" swimtime="00:01:37.10" />
                    <SPLIT distance="200" swimtime="00:01:52.71" />
                    <SPLIT distance="225" swimtime="00:02:03.51" />
                    <SPLIT distance="250" swimtime="00:02:16.51" />
                    <SPLIT distance="275" swimtime="00:02:30.44" />
                    <SPLIT distance="300" swimtime="00:02:44.85" />
                    <SPLIT distance="325" swimtime="00:02:55.65" />
                    <SPLIT distance="350" swimtime="00:03:08.54" />
                    <SPLIT distance="375" swimtime="00:03:21.66" />
                    <SPLIT distance="400" swimtime="00:03:34.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="122443" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="156135" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="197192" reactiontime="+33" />
                    <RELAYPOSITION number="4" athleteid="150083" reactiontime="+13" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="Turkey">
              <RESULTS>
                <RESULT eventid="11" place="19" lane="3" heat="4" swimtime="00:01:44.49" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:24.64" />
                    <SPLIT distance="75" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:00:50.35" />
                    <SPLIT distance="125" swimtime="00:01:02.85" />
                    <SPLIT distance="150" swimtime="00:01:17.69" />
                    <SPLIT distance="175" swimtime="00:01:30.50" />
                    <SPLIT distance="200" swimtime="00:01:44.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="122443" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="110514" reactiontime="+5" />
                    <RELAYPOSITION number="3" athleteid="110602" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="170682" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Turkey">
              <RESULTS>
                <RESULT eventid="35" place="13" lane="3" heat="3" swimtime="00:01:35.23" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.91" />
                    <SPLIT distance="50" swimtime="00:00:24.42" />
                    <SPLIT distance="75" swimtime="00:00:36.45" />
                    <SPLIT distance="100" swimtime="00:00:50.81" />
                    <SPLIT distance="125" swimtime="00:01:01.09" />
                    <SPLIT distance="150" swimtime="00:01:13.93" />
                    <SPLIT distance="175" swimtime="00:01:23.96" />
                    <SPLIT distance="200" swimtime="00:01:35.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="122443" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="156135" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="150083" reactiontime="+3" />
                    <RELAYPOSITION number="4" athleteid="110514" reactiontime="+16" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Utd Arab Emirates" shortname="UAE" code="UAE" nation="UAE" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="129079" lastname="ALHAMMADI" firstname="Omar Mohammed Ahmed Mohammed" gender="M" birthdate="1993-04-18">
              <ENTRIES>
                <ENTRY entrytime="00:01:05.48" eventid="16" heat="2" lane="8">
                  <MEETINFO date="2021-10-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.05" eventid="41" heat="2" lane="4">
                  <MEETINFO date="2021-10-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="54" lane="8" heat="2" heatid="20016" swimtime="00:01:04.57" reactiontime="+74" points="627">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                    <SPLIT distance="75" swimtime="00:00:47.08" />
                    <SPLIT distance="100" swimtime="00:01:04.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="52" lane="4" heat="2" heatid="20041" swimtime="00:00:29.96" reactiontime="+69" points="577">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.86" />
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="164374" lastname="SABT" firstname="Salem" gender="M" birthdate="2005-05-19">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.15" eventid="39" heat="2" lane="3">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:52.46" eventid="14" heat="4" lane="8">
                  <MEETINFO date="2022-08-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="44" lane="3" heat="2" heatid="20039" swimtime="00:00:55.95" reactiontime="+67" points="622">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.83" />
                    <SPLIT distance="50" swimtime="00:00:25.85" />
                    <SPLIT distance="75" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:00:55.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="55" lane="8" heat="4" heatid="40014" swimtime="00:00:50.58" reactiontime="+69" points="696">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.46" />
                    <SPLIT distance="50" swimtime="00:00:24.17" />
                    <SPLIT distance="75" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213783" lastname="ALSHEHHI" firstname="Mahra" gender="F" birthdate="2006-07-12">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="13" heat="1" lane="3" />
                <ENTRY entrytime="NT" eventid="30" heat="1" lane="2" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="-1" lane="3" heat="1" heatid="10013" swimtime="NT" status="DNS" />
                <RESULT eventid="30" place="-1" lane="2" heat="1" heatid="10030" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213782" lastname="ALSHEHHI" firstname="Maha" gender="F" birthdate="2006-07-12">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="43" heat="1" lane="8" />
                <ENTRY entrytime="NT" eventid="1" heat="1" lane="1" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="43" place="-1" lane="8" heat="1" heatid="10043" swimtime="NT" status="DNS" />
                <RESULT eventid="1" place="-1" lane="1" heat="1" heatid="10001" swimtime="NT" status="DNS" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Uganda" shortname="UGA" code="UGA" nation="UGA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="153516" lastname="SSENGONZI" firstname="Jesse Ssuubi" gender="M" birthdate="2002-08-27">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.64" eventid="39" heat="4" lane="8">
                  <MEETINFO date="2021-12-17" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.15" eventid="5" heat="4" lane="5">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="29" lane="8" heat="4" heatid="40039" swimtime="00:00:51.90" reactiontime="+62" points="780">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.91" />
                    <SPLIT distance="50" swimtime="00:00:24.02" />
                    <SPLIT distance="75" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:00:51.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="48" lane="5" heat="4" heatid="40005" swimtime="00:00:23.79" reactiontime="+64" points="764">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.89" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="211075" lastname="NALUWOZA" firstname="Tara Ann Mary" gender="F" birthdate="2008-08-05">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="38" heat="1" lane="1" />
                <ENTRY entrytime="00:00:28.97" eventid="4" heat="3" lane="1">
                  <MEETINFO date="2022-09-01" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="38" place="29" lane="1" heat="1" heatid="10038" swimtime="00:01:05.28" reactiontime="+71" points="584">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="75" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="30" lane="1" heat="3" heatid="30004" swimtime="00:00:27.71" reactiontime="+74" points="681">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.81" />
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="153511" lastname="NAMUTEBI" firstname="Kirabo" gender="F" birthdate="2005-02-08">
              <ENTRIES>
                <ENTRY entrytime="00:00:33.25" eventid="40" heat="3" lane="5">
                  <MEETINFO date="2021-10-30" />
                </ENTRY>
                <ENTRY entrytime="00:00:25.84" eventid="30" heat="4" lane="5">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="40" place="29" lane="5" heat="3" heatid="30040" swimtime="00:00:32.47" reactiontime="+64" points="680">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.71" />
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="34" lane="5" heat="4" heatid="40030" swimtime="00:00:26.15" reactiontime="+64" points="674">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.58" />
                    <SPLIT distance="50" swimtime="00:00:26.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Ukraine" shortname="UKR" code="UKR" nation="UKR" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="197925" lastname="LISOVETS" firstname="Volodymyr" gender="M" birthdate="2004-05-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.25" eventid="16" heat="4" lane="2">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:27.34" eventid="41" heat="5" lane="5">
                  <MEETINFO date="2022-08-15" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="35" lane="2" heat="4" heatid="40016" swimtime="00:00:59.55" reactiontime="+67" points="799">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.63" />
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="75" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:00:59.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="26" lane="5" heat="5" heatid="50041" swimtime="00:00:27.04" reactiontime="+67" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.31" />
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183260" lastname="LINNYK" firstname="Illia" gender="M" birthdate="2001-03-14">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.10" eventid="14" heat="8" lane="8">
                  <MEETINFO date="2022-10-22" />
                </ENTRY>
                <ENTRY entrytime="00:01:46.88" eventid="44" heat="3" lane="8">
                  <MEETINFO date="2021-10-22" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:22.18" eventid="31" heat="6" lane="4">
                  <MEETINFO date="2022-08-16" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="39" lane="8" heat="8" heatid="80014" swimtime="00:00:47.99" reactiontime="+68" points="815">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.61" />
                    <SPLIT distance="50" swimtime="00:00:22.75" />
                    <SPLIT distance="75" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="34" lane="8" heat="3" heatid="30044" swimtime="00:01:47.72" reactiontime="+68" points="785">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                    <SPLIT distance="75" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:00:52.14" />
                    <SPLIT distance="125" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:19.88" />
                    <SPLIT distance="175" swimtime="00:01:34.13" />
                    <SPLIT distance="200" swimtime="00:01:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="41" lane="4" heat="6" heatid="60031" swimtime="00:00:21.73" reactiontime="+66" points="798">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.53" />
                    <SPLIT distance="50" swimtime="00:00:21.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="102652" lastname="GOVOROV" firstname="Andrii" gender="M" birthdate="1992-04-10">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.18" eventid="5" heat="7" lane="8">
                  <MEETINFO date="2022-08-12" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="5" place="29" lane="8" heat="7" heatid="70005" swimtime="00:00:22.92" reactiontime="+61" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:22.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="182982" lastname="BUKHOV" firstname="Vladyslav" gender="M" birthdate="2002-07-05">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.16" eventid="31" heat="10" lane="6">
                  <MEETINFO date="2021-09-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="10" lane="6" heat="10" heatid="100031" swimtime="00:00:21.13" reactiontime="+70" points="868">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="231" place="14" lane="2" heat="2" heatid="20231" swimtime="00:00:21.29" reactiontime="+70" points="849">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.24" />
                    <SPLIT distance="50" swimtime="00:00:21.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197926" lastname="ZHELTIAKOV" firstname="Oleksandr" gender="M" birthdate="2005-11-15" />
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Ukraine">
              <RESULTS>
                <RESULT eventid="48" place="16" lane="1" heat="3" swimtime="00:03:37.84" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.56" />
                    <SPLIT distance="50" swimtime="00:00:26.38" />
                    <SPLIT distance="75" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:00:54.47" />
                    <SPLIT distance="125" swimtime="00:01:07.03" />
                    <SPLIT distance="150" swimtime="00:01:22.46" />
                    <SPLIT distance="175" swimtime="00:01:38.40" />
                    <SPLIT distance="200" swimtime="00:01:55.12" />
                    <SPLIT distance="225" swimtime="00:02:05.77" />
                    <SPLIT distance="250" swimtime="00:02:19.41" />
                    <SPLIT distance="275" swimtime="00:02:33.95" />
                    <SPLIT distance="300" swimtime="00:02:49.62" />
                    <SPLIT distance="325" swimtime="00:03:00.14" />
                    <SPLIT distance="350" swimtime="00:03:12.25" />
                    <SPLIT distance="375" swimtime="00:03:25.24" />
                    <SPLIT distance="400" swimtime="00:03:37.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197926" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="197925" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="102652" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="183260" reactiontime="+43" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Ukraine">
              <RESULTS>
                <RESULT eventid="126" place="7" lane="8" heat="1" swimtime="00:01:26.11" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.41" />
                    <SPLIT distance="50" swimtime="00:00:21.78" />
                    <SPLIT distance="75" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:00:42.90" />
                    <SPLIT distance="125" swimtime="00:00:52.59" />
                    <SPLIT distance="150" swimtime="00:01:03.37" />
                    <SPLIT distance="175" swimtime="00:01:13.98" />
                    <SPLIT distance="200" swimtime="00:01:26.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="102652" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="183260" reactiontime="+27" />
                    <RELAYPOSITION number="3" athleteid="182982" reactiontime="+9" />
                    <RELAYPOSITION number="4" athleteid="197926" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="8" lane="2" heat="2" swimtime="00:01:26.53" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.36" />
                    <SPLIT distance="50" swimtime="00:00:21.70" />
                    <SPLIT distance="75" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:00:42.67" />
                    <SPLIT distance="125" swimtime="00:00:52.56" />
                    <SPLIT distance="150" swimtime="00:01:03.61" />
                    <SPLIT distance="175" swimtime="00:01:14.27" />
                    <SPLIT distance="200" swimtime="00:01:26.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="102652" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="183260" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="182982" reactiontime="+11" />
                    <RELAYPOSITION number="4" athleteid="197926" reactiontime="+33" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="Ukraine">
              <RESULTS>
                <RESULT eventid="35" place="9" lane="3" heat="2" swimtime="00:01:34.35" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:24.25" />
                    <SPLIT distance="75" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:00:50.69" />
                    <SPLIT distance="125" swimtime="00:01:00.81" />
                    <SPLIT distance="150" swimtime="00:01:13.45" />
                    <SPLIT distance="175" swimtime="00:01:23.39" />
                    <SPLIT distance="200" swimtime="00:01:34.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197926" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="197925" reactiontime="+23" />
                    <RELAYPOSITION number="3" athleteid="102652" reactiontime="+19" />
                    <RELAYPOSITION number="4" athleteid="182982" reactiontime="+14" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Uruguay" shortname="URU" code="URU" nation="URU" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="123478" lastname="CHIANCONE" firstname="Pedro" gender="M" birthdate="1997-07-20">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.18" eventid="14" heat="6" lane="2">
                  <MEETINFO date="2021-10-28" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="52" lane="2" heat="6" heatid="60014" swimtime="00:00:50.28" reactiontime="+63" points="709">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.36" />
                    <SPLIT distance="50" swimtime="00:00:23.86" />
                    <SPLIT distance="75" swimtime="00:00:36.97" />
                    <SPLIT distance="100" swimtime="00:00:50.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="100884" lastname="MELCONIAN" firstname="Martin" gender="M" birthdate="1990-01-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:27.93" eventid="41" heat="4" lane="5">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="41" place="41" lane="5" heat="4" heatid="40041" swimtime="00:00:27.79" reactiontime="+62" points="723">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="123670" lastname="AUNCHAYNA" firstname="Aabril" gender="F" birthdate="1999-04-08">
              <ENTRIES>
                <ENTRY entrytime="00:01:06.87" eventid="2" heat="2" lane="8">
                  <MEETINFO date="2022-05-07" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.20" eventid="18" heat="3" lane="7">
                  <MEETINFO date="2022-03-23" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="32" lane="8" heat="2" heatid="20002" swimtime="00:01:01.07" reactiontime="+57" points="726">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.81" />
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="75" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:01.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="29" lane="7" heat="3" heatid="30018" swimtime="00:00:28.06" reactiontime="+56" points="730">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.80" />
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="169845" lastname="FRANK" firstname="Nicole" gender="F" birthdate="2003-09-08">
              <ENTRIES>
                <ENTRY entrytime="00:02:33.36" eventid="28" heat="1" lane="5">
                  <MEETINFO date="2021-11-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="28" place="24" lane="5" heat="1" heatid="10028" swimtime="00:02:26.44" reactiontime="+65" points="776">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.15" />
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="75" swimtime="00:00:51.17" />
                    <SPLIT distance="100" swimtime="00:01:09.49" />
                    <SPLIT distance="125" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:01:47.35" />
                    <SPLIT distance="175" swimtime="00:02:06.94" />
                    <SPLIT distance="200" swimtime="00:02:26.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="United States" shortname="USA" code="USA" nation="USA" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="105644" lastname="MURPHY" firstname="Ryan" gender="M" birthdate="1995-07-02">
              <ENTRIES>
                <ENTRY entrytime="00:00:49.44" eventid="3" heat="4" lane="4">
                  <MEETINFO date="2021-11-13" />
                </ENTRY>
                <ENTRY entrytime="00:01:48.10" eventid="46" heat="4" lane="4">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:22.53" eventid="19" heat="6" lane="4">
                  <MEETINFO date="2021-11-25" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="103" place="1" lane="4" heat="1" heatid="10103" swimtime="00:00:48.50" reactiontime="+50" points="989">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.37" />
                    <SPLIT distance="50" swimtime="00:00:23.40" />
                    <SPLIT distance="75" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:00:48.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="3" place="1" lane="4" heat="4" heatid="40003" swimtime="00:00:49.34" reactiontime="+50" points="939">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.50" />
                    <SPLIT distance="50" swimtime="00:00:23.66" />
                    <SPLIT distance="75" swimtime="00:00:36.47" />
                    <SPLIT distance="100" swimtime="00:00:49.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="203" place="1" lane="4" heat="2" heatid="20203" swimtime="00:00:49.17" reactiontime="+49" points="949">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                    <SPLIT distance="75" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:00:49.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="146" place="1" lane="3" heat="1" heatid="10146" swimtime="00:01:47.41" reactiontime="+52" points="951">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.84" />
                    <SPLIT distance="50" swimtime="00:00:25.09" />
                    <SPLIT distance="75" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:00:52.22" />
                    <SPLIT distance="125" swimtime="00:01:05.82" />
                    <SPLIT distance="150" swimtime="00:01:19.50" />
                    <SPLIT distance="175" swimtime="00:01:33.24" />
                    <SPLIT distance="200" swimtime="00:01:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="3" lane="4" heat="4" heatid="40046" swimtime="00:01:49.71" reactiontime="+55" points="892">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.19" />
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                    <SPLIT distance="75" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:00:53.68" />
                    <SPLIT distance="125" swimtime="00:01:07.74" />
                    <SPLIT distance="150" swimtime="00:01:21.85" />
                    <SPLIT distance="175" swimtime="00:01:36.08" />
                    <SPLIT distance="200" swimtime="00:01:49.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="119" place="1" lane="5" heat="1" heatid="10119" swimtime="00:00:22.64" reactiontime="+51" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.12" />
                    <SPLIT distance="50" swimtime="00:00:22.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="10" lane="4" heat="6" heatid="60019" swimtime="00:00:23.22" reactiontime="+51" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.54" />
                    <SPLIT distance="50" swimtime="00:00:23.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="2" lane="2" heat="1" heatid="10219" swimtime="00:00:22.74" reactiontime="+52" points="932">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.09" />
                    <SPLIT distance="50" swimtime="00:00:22.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183481" lastname="ARMSTRONG" firstname="Hunter" gender="M" birthdate="2001-01-24">
              <ENTRIES>
                <ENTRY entrytime="00:00:51.98" eventid="3" heat="4" lane="8">
                  <MEETINFO date="2022-06-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:48.25" eventid="14" heat="7" lane="4">
                  <MEETINFO date="2022-04-26" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:23.70" eventid="19" heat="6" lane="8">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="3" place="17" lane="8" heat="4" heatid="40003" swimtime="00:00:50.93" reactiontime="+64" points="854">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.94" />
                    <SPLIT distance="50" swimtime="00:00:24.77" />
                    <SPLIT distance="75" swimtime="00:00:37.85" />
                    <SPLIT distance="100" swimtime="00:00:50.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="14" place="19" lane="4" heat="7" heatid="70014" swimtime="00:00:47.11" reactiontime="+64" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.72" />
                    <SPLIT distance="50" swimtime="00:00:22.80" />
                    <SPLIT distance="75" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="19" place="8" lane="8" heat="6" heatid="60019" swimtime="00:00:23.18" reactiontime="+59" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.32" />
                    <SPLIT distance="50" swimtime="00:00:23.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="219" place="8" lane="2" heat="2" heatid="20219" swimtime="00:00:23.05" reactiontime="+58" points="895">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.25" />
                    <SPLIT distance="50" swimtime="00:00:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="419" place="9" lane="5" heat="1" heatid="10419" swimtime="00:00:23.30" reactiontime="+57" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:23.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105614" lastname="FINK" firstname="Nic" gender="M" birthdate="1993-07-03">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.56" eventid="16" heat="8" lane="4">
                  <MEETINFO date="2021-12-04" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.28" eventid="29" heat="5" lane="5">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="00:00:25.53" eventid="41" heat="7" lane="4">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="116" place="1" lane="5" heat="1" heatid="10116" swimtime="00:00:55.88" reactiontime="+71" points="968">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:26.04" />
                    <SPLIT distance="75" swimtime="00:00:40.72" />
                    <SPLIT distance="100" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="16" place="5" lane="4" heat="8" heatid="80016" swimtime="00:00:57.02" reactiontime="+72" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.13" />
                    <SPLIT distance="50" swimtime="00:00:26.68" />
                    <SPLIT distance="75" swimtime="00:00:41.63" />
                    <SPLIT distance="100" swimtime="00:00:57.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="216" place="2" lane="3" heat="2" heatid="20216" swimtime="00:00:56.25" reactiontime="+71" points="949">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                    <SPLIT distance="50" swimtime="00:00:26.29" />
                    <SPLIT distance="75" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:00:56.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="129" place="2" lane="5" heat="1" heatid="10129" swimtime="00:02:01.60" reactiontime="+71" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.43" />
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                    <SPLIT distance="75" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:00:59.04" />
                    <SPLIT distance="125" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:30.23" />
                    <SPLIT distance="175" swimtime="00:01:45.63" />
                    <SPLIT distance="200" swimtime="00:02:01.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="29" place="2" lane="5" heat="5" heatid="50029" swimtime="00:02:02.75" reactiontime="+72" points="938">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.68" />
                    <SPLIT distance="50" swimtime="00:00:28.03" />
                    <SPLIT distance="75" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:00:59.95" />
                    <SPLIT distance="125" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:31.70" />
                    <SPLIT distance="175" swimtime="00:01:47.19" />
                    <SPLIT distance="200" swimtime="00:02:02.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="1" lane="5" heat="1" heatid="10141" swimtime="00:00:25.38" reactiontime="+71" points="950">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="4" lane="4" heat="7" heatid="70041" swimtime="00:00:26.07" reactiontime="+70" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="2" lane="5" heat="1" heatid="10241" swimtime="00:00:25.64" reactiontime="+69" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                    <SPLIT distance="50" swimtime="00:00:25.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124916" lastname="ANDREW" firstname="Michael" gender="M" birthdate="1999-04-18">
              <ENTRIES>
                <ENTRY entrytime="00:00:57.54" eventid="16" heat="8" lane="1">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:00:50.88" eventid="39" heat="5" lane="4">
                  <MEETINFO date="2022-04-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:26.32" eventid="41" heat="7" lane="2">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:00:22.79" eventid="5" heat="7" lane="4">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.41" eventid="31" heat="8" lane="5">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:51.22" eventid="23" heat="4" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="25" lane="1" heat="8" heatid="80016" swimtime="00:00:58.22" reactiontime="+67" points="856">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.88" />
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                    <SPLIT distance="75" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:00:58.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="39" place="30" lane="4" heat="5" heatid="50039" swimtime="00:00:51.93" reactiontime="+75" points="778">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.60" />
                    <SPLIT distance="50" swimtime="00:00:23.57" />
                    <SPLIT distance="75" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:00:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="141" place="5" lane="2" heat="1" heatid="10141" swimtime="00:00:25.92" reactiontime="+70" points="891">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.52" />
                    <SPLIT distance="50" swimtime="00:00:25.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="41" place="8" lane="2" heat="7" heatid="70041" swimtime="00:00:26.17" reactiontime="+67" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                    <SPLIT distance="50" swimtime="00:00:26.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="241" place="5" lane="6" heat="1" heatid="10241" swimtime="00:00:25.81" reactiontime="+66" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.55" />
                    <SPLIT distance="50" swimtime="00:00:25.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="10" lane="4" heat="7" heatid="70005" swimtime="00:00:22.34" reactiontime="+67" points="922">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.98" />
                    <SPLIT distance="50" swimtime="00:00:22.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="205" place="14" lane="2" heat="1" heatid="10205" swimtime="00:00:22.47" reactiontime="+67" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.04" />
                    <SPLIT distance="50" swimtime="00:00:22.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="8" lane="5" heat="8" heatid="80031" swimtime="00:00:21.02" reactiontime="+68" points="882">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.09" />
                    <SPLIT distance="50" swimtime="00:00:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="5" lane="4" heat="1" heatid="10123" swimtime="00:00:51.47" reactiontime="+66" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.19" />
                    <SPLIT distance="50" swimtime="00:00:23.12" />
                    <SPLIT distance="75" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:00:51.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="7" lane="4" heat="4" heatid="40023" swimtime="00:00:52.21" reactiontime="+68" points="840">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.40" />
                    <SPLIT distance="50" swimtime="00:00:23.42" />
                    <SPLIT distance="75" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:00:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="1" lane="6" heat="2" heatid="20223" swimtime="00:00:51.40" reactiontime="+67" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.21" />
                    <SPLIT distance="50" swimtime="00:00:23.22" />
                    <SPLIT distance="75" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:00:51.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197510" lastname="CASAS" firstname="Shaine" gender="M" birthdate="1999-12-25">
              <ENTRIES>
                <ENTRY entrytime="00:00:50.40" eventid="39" heat="7" lane="1">
                  <MEETINFO date="2022-07-28" />
                </ENTRY>
                <ENTRY entrytime="00:01:48.40" eventid="46" heat="3" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="00:01:50.37" eventid="7" heat="5" lane="4">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:51.03" eventid="23" heat="5" lane="4">
                  <MEETINFO date="2022-10-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="11" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="-1" lane="1" heat="7" heatid="70039" swimtime="NT" status="DNS" />
                <RESULT eventid="146" place="2" lane="4" heat="1" heatid="10146" swimtime="00:01:48.01" reactiontime="+51" points="935">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.86" />
                    <SPLIT distance="50" swimtime="00:00:25.02" />
                    <SPLIT distance="75" swimtime="00:00:38.64" />
                    <SPLIT distance="100" swimtime="00:00:52.57" />
                    <SPLIT distance="125" swimtime="00:01:06.39" />
                    <SPLIT distance="150" swimtime="00:01:20.24" />
                    <SPLIT distance="175" swimtime="00:01:34.25" />
                    <SPLIT distance="200" swimtime="00:01:48.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="46" place="1" lane="4" heat="3" heatid="30046" swimtime="00:01:49.46" reactiontime="+52" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.90" />
                    <SPLIT distance="50" swimtime="00:00:25.04" />
                    <SPLIT distance="75" swimtime="00:00:38.92" />
                    <SPLIT distance="100" swimtime="00:00:52.80" />
                    <SPLIT distance="125" swimtime="00:01:06.92" />
                    <SPLIT distance="150" swimtime="00:01:20.96" />
                    <SPLIT distance="175" swimtime="00:01:35.36" />
                    <SPLIT distance="200" swimtime="00:01:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="107" place="4" lane="2" heat="1" heatid="10107" swimtime="00:01:51.31" reactiontime="+62" points="955">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.65" />
                    <SPLIT distance="50" swimtime="00:00:23.57" />
                    <SPLIT distance="75" swimtime="00:00:37.86" />
                    <SPLIT distance="100" swimtime="00:00:51.06" />
                    <SPLIT distance="125" swimtime="00:01:07.06" />
                    <SPLIT distance="150" swimtime="00:01:23.48" />
                    <SPLIT distance="175" swimtime="00:01:37.96" />
                    <SPLIT distance="200" swimtime="00:01:51.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="4" lane="4" heat="5" heatid="50007" swimtime="00:01:52.52" reactiontime="+61" points="924">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:23.79" />
                    <SPLIT distance="75" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:00:52.02" />
                    <SPLIT distance="125" swimtime="00:01:08.15" />
                    <SPLIT distance="150" swimtime="00:01:24.77" />
                    <SPLIT distance="175" swimtime="00:01:39.33" />
                    <SPLIT distance="200" swimtime="00:01:52.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="123" place="4" lane="5" heat="1" heatid="10123" swimtime="00:00:51.36" reactiontime="+59" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.43" />
                    <SPLIT distance="50" swimtime="00:00:23.08" />
                    <SPLIT distance="75" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:00:51.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="23" place="3" lane="4" heat="5" heatid="50023" swimtime="00:00:51.96" reactiontime="+62" points="853">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.52" />
                    <SPLIT distance="50" swimtime="00:00:23.27" />
                    <SPLIT distance="75" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:00:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="223" place="2" lane="5" heat="2" heatid="20223" swimtime="00:00:51.42" reactiontime="+61" points="880">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.35" />
                    <SPLIT distance="50" swimtime="00:00:22.95" />
                    <SPLIT distance="75" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:00:51.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="145806" lastname="KIBLER" firstname="Drew" gender="M" birthdate="2000-03-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:46.82" eventid="14" heat="9" lane="2">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:41.93" eventid="44" heat="6" lane="3">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="26" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="17" lane="2" heat="9" heatid="90014" swimtime="00:00:47.05" reactiontime="+63" points="865">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.68" />
                    <SPLIT distance="50" swimtime="00:00:22.64" />
                    <SPLIT distance="75" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:00:47.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="144" place="4" lane="6" heat="1" heatid="10144" swimtime="00:01:41.44" reactiontime="+63" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.18" />
                    <SPLIT distance="50" swimtime="00:00:23.68" />
                    <SPLIT distance="75" swimtime="00:00:36.39" />
                    <SPLIT distance="100" swimtime="00:00:49.38" />
                    <SPLIT distance="125" swimtime="00:01:02.40" />
                    <SPLIT distance="150" swimtime="00:01:15.56" />
                    <SPLIT distance="175" swimtime="00:01:28.69" />
                    <SPLIT distance="200" swimtime="00:01:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="44" place="4" lane="3" heat="6" heatid="60044" swimtime="00:01:41.88" reactiontime="+63" points="927">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.11" />
                    <SPLIT distance="50" swimtime="00:00:23.77" />
                    <SPLIT distance="75" swimtime="00:00:36.65" />
                    <SPLIT distance="100" swimtime="00:00:49.50" />
                    <SPLIT distance="125" swimtime="00:01:02.40" />
                    <SPLIT distance="150" swimtime="00:01:15.56" />
                    <SPLIT distance="175" swimtime="00:01:28.89" />
                    <SPLIT distance="200" swimtime="00:01:41.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202563" lastname="CLARK" firstname="Charlie" gender="M" birthdate="2002-06-17">
              <ENTRIES>
                <ENTRY entrytime="00:14:51.78" eventid="10" heat="2" lane="1">
                  <MEETINFO date="2022-04-26" />
                </ENTRY>
                <ENTRY entrytime="00:07:50.07" eventid="42" heat="2" lane="7">
                  <MEETINFO date="2022-04-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="7" lane="1" heat="2" heatid="20010" swimtime="00:14:33.93" reactiontime="+66" points="909">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:26.99" />
                    <SPLIT distance="75" swimtime="00:00:41.40" />
                    <SPLIT distance="100" swimtime="00:00:55.98" />
                    <SPLIT distance="125" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:25.35" />
                    <SPLIT distance="175" swimtime="00:01:39.90" />
                    <SPLIT distance="200" swimtime="00:01:54.65" />
                    <SPLIT distance="225" swimtime="00:02:09.26" />
                    <SPLIT distance="250" swimtime="00:02:24.02" />
                    <SPLIT distance="275" swimtime="00:02:38.60" />
                    <SPLIT distance="300" swimtime="00:02:53.36" />
                    <SPLIT distance="325" swimtime="00:03:08.02" />
                    <SPLIT distance="350" swimtime="00:03:22.79" />
                    <SPLIT distance="375" swimtime="00:03:37.45" />
                    <SPLIT distance="400" swimtime="00:03:52.34" />
                    <SPLIT distance="425" swimtime="00:04:06.96" />
                    <SPLIT distance="450" swimtime="00:04:21.75" />
                    <SPLIT distance="475" swimtime="00:04:36.28" />
                    <SPLIT distance="500" swimtime="00:04:50.98" />
                    <SPLIT distance="525" swimtime="00:05:05.56" />
                    <SPLIT distance="550" swimtime="00:05:20.41" />
                    <SPLIT distance="575" swimtime="00:05:35.05" />
                    <SPLIT distance="600" swimtime="00:05:49.82" />
                    <SPLIT distance="625" swimtime="00:06:04.44" />
                    <SPLIT distance="650" swimtime="00:06:19.19" />
                    <SPLIT distance="675" swimtime="00:06:33.80" />
                    <SPLIT distance="700" swimtime="00:06:48.45" />
                    <SPLIT distance="725" swimtime="00:07:03.08" />
                    <SPLIT distance="750" swimtime="00:07:17.69" />
                    <SPLIT distance="775" swimtime="00:07:32.29" />
                    <SPLIT distance="800" swimtime="00:07:46.91" />
                    <SPLIT distance="825" swimtime="00:08:01.48" />
                    <SPLIT distance="850" swimtime="00:08:16.08" />
                    <SPLIT distance="875" swimtime="00:08:30.63" />
                    <SPLIT distance="900" swimtime="00:08:45.27" />
                    <SPLIT distance="925" swimtime="00:08:59.82" />
                    <SPLIT distance="950" swimtime="00:09:14.45" />
                    <SPLIT distance="975" swimtime="00:09:29.04" />
                    <SPLIT distance="1000" swimtime="00:09:43.66" />
                    <SPLIT distance="1025" swimtime="00:09:58.29" />
                    <SPLIT distance="1050" swimtime="00:10:12.91" />
                    <SPLIT distance="1075" swimtime="00:10:27.46" />
                    <SPLIT distance="1100" swimtime="00:10:42.04" />
                    <SPLIT distance="1125" swimtime="00:10:56.59" />
                    <SPLIT distance="1150" swimtime="00:11:11.23" />
                    <SPLIT distance="1175" swimtime="00:11:25.87" />
                    <SPLIT distance="1200" swimtime="00:11:40.57" />
                    <SPLIT distance="1225" swimtime="00:11:55.17" />
                    <SPLIT distance="1250" swimtime="00:12:09.89" />
                    <SPLIT distance="1275" swimtime="00:12:24.51" />
                    <SPLIT distance="1300" swimtime="00:12:39.17" />
                    <SPLIT distance="1325" swimtime="00:12:53.76" />
                    <SPLIT distance="1350" swimtime="00:13:08.42" />
                    <SPLIT distance="1375" swimtime="00:13:22.98" />
                    <SPLIT distance="1400" swimtime="00:13:37.47" />
                    <SPLIT distance="1425" swimtime="00:13:51.72" />
                    <SPLIT distance="1450" swimtime="00:14:06.13" />
                    <SPLIT distance="1475" swimtime="00:14:20.30" />
                    <SPLIT distance="1500" swimtime="00:14:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="8" lane="7" heat="2" heatid="20042" swimtime="00:07:37.54" reactiontime="+67" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.36" />
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                    <SPLIT distance="75" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:00:55.55" />
                    <SPLIT distance="125" swimtime="00:01:10.05" />
                    <SPLIT distance="150" swimtime="00:01:24.70" />
                    <SPLIT distance="175" swimtime="00:01:39.23" />
                    <SPLIT distance="200" swimtime="00:01:53.83" />
                    <SPLIT distance="225" swimtime="00:02:08.27" />
                    <SPLIT distance="250" swimtime="00:02:22.80" />
                    <SPLIT distance="275" swimtime="00:02:37.30" />
                    <SPLIT distance="300" swimtime="00:02:51.75" />
                    <SPLIT distance="325" swimtime="00:03:06.15" />
                    <SPLIT distance="350" swimtime="00:03:20.65" />
                    <SPLIT distance="375" swimtime="00:03:35.05" />
                    <SPLIT distance="400" swimtime="00:03:49.45" />
                    <SPLIT distance="425" swimtime="00:04:03.70" />
                    <SPLIT distance="450" swimtime="00:04:18.00" />
                    <SPLIT distance="475" swimtime="00:04:32.40" />
                    <SPLIT distance="500" swimtime="00:04:46.70" />
                    <SPLIT distance="525" swimtime="00:05:00.86" />
                    <SPLIT distance="550" swimtime="00:05:15.10" />
                    <SPLIT distance="575" swimtime="00:05:29.39" />
                    <SPLIT distance="600" swimtime="00:05:43.59" />
                    <SPLIT distance="625" swimtime="00:05:57.78" />
                    <SPLIT distance="650" swimtime="00:06:11.92" />
                    <SPLIT distance="675" swimtime="00:06:26.27" />
                    <SPLIT distance="700" swimtime="00:06:40.59" />
                    <SPLIT distance="725" swimtime="00:06:54.90" />
                    <SPLIT distance="750" swimtime="00:07:09.41" />
                    <SPLIT distance="775" swimtime="00:07:23.75" />
                    <SPLIT distance="800" swimtime="00:07:37.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214520" lastname="JOHNSTON" firstname="David" gender="M" birthdate="2001-10-28">
              <ENTRIES>
                <ENTRY entrytime="00:14:22.77" eventid="10" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
                <ENTRY entrytime="00:07:30.41" eventid="42" heat="0" lane="2147483647">
                  <MEETINFO date="2022-08-24" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="110" place="8" lane="5" heat="5" heatid="30110" swimtime="00:14:35.27" reactiontime="+73" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                    <SPLIT distance="75" swimtime="00:00:40.86" />
                    <SPLIT distance="100" swimtime="00:00:55.05" />
                    <SPLIT distance="125" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:23.83" />
                    <SPLIT distance="175" swimtime="00:01:38.32" />
                    <SPLIT distance="200" swimtime="00:01:52.83" />
                    <SPLIT distance="225" swimtime="00:02:07.38" />
                    <SPLIT distance="250" swimtime="00:02:22.01" />
                    <SPLIT distance="275" swimtime="00:02:36.69" />
                    <SPLIT distance="300" swimtime="00:02:51.20" />
                    <SPLIT distance="325" swimtime="00:03:05.81" />
                    <SPLIT distance="350" swimtime="00:03:20.23" />
                    <SPLIT distance="375" swimtime="00:03:34.89" />
                    <SPLIT distance="400" swimtime="00:03:49.42" />
                    <SPLIT distance="425" swimtime="00:04:04.12" />
                    <SPLIT distance="450" swimtime="00:04:18.72" />
                    <SPLIT distance="475" swimtime="00:04:33.41" />
                    <SPLIT distance="500" swimtime="00:04:47.96" />
                    <SPLIT distance="525" swimtime="00:05:02.64" />
                    <SPLIT distance="550" swimtime="00:05:17.19" />
                    <SPLIT distance="575" swimtime="00:05:31.90" />
                    <SPLIT distance="600" swimtime="00:05:46.43" />
                    <SPLIT distance="625" swimtime="00:06:01.20" />
                    <SPLIT distance="650" swimtime="00:06:15.70" />
                    <SPLIT distance="675" swimtime="00:06:30.46" />
                    <SPLIT distance="700" swimtime="00:06:45.02" />
                    <SPLIT distance="725" swimtime="00:06:59.76" />
                    <SPLIT distance="750" swimtime="00:07:14.28" />
                    <SPLIT distance="775" swimtime="00:07:28.90" />
                    <SPLIT distance="800" swimtime="00:07:43.40" />
                    <SPLIT distance="825" swimtime="00:07:58.00" />
                    <SPLIT distance="850" swimtime="00:08:12.48" />
                    <SPLIT distance="875" swimtime="00:08:27.15" />
                    <SPLIT distance="900" swimtime="00:08:41.73" />
                    <SPLIT distance="925" swimtime="00:08:56.45" />
                    <SPLIT distance="950" swimtime="00:09:10.93" />
                    <SPLIT distance="975" swimtime="00:09:25.67" />
                    <SPLIT distance="1000" swimtime="00:09:40.23" />
                    <SPLIT distance="1025" swimtime="00:09:54.93" />
                    <SPLIT distance="1050" swimtime="00:10:09.48" />
                    <SPLIT distance="1075" swimtime="00:10:24.08" />
                    <SPLIT distance="1100" swimtime="00:10:38.72" />
                    <SPLIT distance="1125" swimtime="00:10:53.59" />
                    <SPLIT distance="1150" swimtime="00:11:08.20" />
                    <SPLIT distance="1175" swimtime="00:11:23.02" />
                    <SPLIT distance="1200" swimtime="00:11:37.72" />
                    <SPLIT distance="1225" swimtime="00:11:52.61" />
                    <SPLIT distance="1250" swimtime="00:12:07.32" />
                    <SPLIT distance="1275" swimtime="00:12:22.23" />
                    <SPLIT distance="1300" swimtime="00:12:36.91" />
                    <SPLIT distance="1325" swimtime="00:12:51.88" />
                    <SPLIT distance="1350" swimtime="00:13:06.86" />
                    <SPLIT distance="1375" swimtime="00:13:21.84" />
                    <SPLIT distance="1400" swimtime="00:13:36.74" />
                    <SPLIT distance="1425" swimtime="00:13:51.69" />
                    <SPLIT distance="1450" swimtime="00:14:06.44" />
                    <SPLIT distance="1475" swimtime="00:14:21.22" />
                    <SPLIT distance="1500" swimtime="00:14:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="142" place="5" lane="5" heat="5" heatid="30142" swimtime="00:07:34.33" reactiontime="+73" points="929">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.39" />
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                    <SPLIT distance="75" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:00:54.32" />
                    <SPLIT distance="125" swimtime="00:01:08.50" />
                    <SPLIT distance="150" swimtime="00:01:22.58" />
                    <SPLIT distance="175" swimtime="00:01:36.95" />
                    <SPLIT distance="200" swimtime="00:01:51.19" />
                    <SPLIT distance="225" swimtime="00:02:05.71" />
                    <SPLIT distance="250" swimtime="00:02:20.05" />
                    <SPLIT distance="275" swimtime="00:02:34.56" />
                    <SPLIT distance="300" swimtime="00:02:48.79" />
                    <SPLIT distance="325" swimtime="00:03:03.20" />
                    <SPLIT distance="350" swimtime="00:03:17.50" />
                    <SPLIT distance="375" swimtime="00:03:31.98" />
                    <SPLIT distance="400" swimtime="00:03:46.32" />
                    <SPLIT distance="425" swimtime="00:04:00.75" />
                    <SPLIT distance="450" swimtime="00:04:14.92" />
                    <SPLIT distance="475" swimtime="00:04:29.25" />
                    <SPLIT distance="500" swimtime="00:04:43.52" />
                    <SPLIT distance="525" swimtime="00:04:57.91" />
                    <SPLIT distance="550" swimtime="00:05:12.26" />
                    <SPLIT distance="575" swimtime="00:05:26.72" />
                    <SPLIT distance="600" swimtime="00:05:40.90" />
                    <SPLIT distance="625" swimtime="00:05:55.17" />
                    <SPLIT distance="650" swimtime="00:06:09.41" />
                    <SPLIT distance="675" swimtime="00:06:23.81" />
                    <SPLIT distance="700" swimtime="00:06:38.03" />
                    <SPLIT distance="725" swimtime="00:06:52.30" />
                    <SPLIT distance="750" swimtime="00:07:06.56" />
                    <SPLIT distance="775" swimtime="00:07:20.79" />
                    <SPLIT distance="800" swimtime="00:07:34.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124840" lastname="SWANSON" firstname="Charlie" gender="M" birthdate="1998-02-20">
              <ENTRIES>
                <ENTRY entrytime="00:02:04.25" eventid="29" heat="3" lane="3">
                  <MEETINFO date="2021-11-11" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="29" place="12" lane="3" heat="3" heatid="30029" swimtime="00:02:05.51" reactiontime="+66" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                    <SPLIT distance="50" swimtime="00:00:28.55" />
                    <SPLIT distance="75" swimtime="00:00:44.07" />
                    <SPLIT distance="100" swimtime="00:01:00.33" />
                    <SPLIT distance="125" swimtime="00:01:16.43" />
                    <SPLIT distance="150" swimtime="00:01:32.73" />
                    <SPLIT distance="175" swimtime="00:01:49.06" />
                    <SPLIT distance="200" swimtime="00:02:05.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124900" lastname="HARTING" firstname="Zach" gender="M" birthdate="1997-08-27">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.74" eventid="21" heat="3" lane="2">
                  <MEETINFO date="2021-11-19" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="21" place="11" lane="2" heat="3" heatid="30021" swimtime="00:01:51.86" reactiontime="+65" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.13" />
                    <SPLIT distance="50" swimtime="00:00:25.00" />
                    <SPLIT distance="75" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:00:53.34" />
                    <SPLIT distance="125" swimtime="00:01:07.69" />
                    <SPLIT distance="150" swimtime="00:01:22.12" />
                    <SPLIT distance="175" swimtime="00:01:36.74" />
                    <SPLIT distance="200" swimtime="00:01:51.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197514" lastname="JULIAN" firstname="Trenton" gender="M" birthdate="1998-12-09">
              <ENTRIES>
                <ENTRY entrytime="00:01:49.69" eventid="21" heat="3" lane="5">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="121" place="7" lane="4" heat="1" heatid="10121" swimtime="00:01:50.94" reactiontime="+63" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.96" />
                    <SPLIT distance="50" swimtime="00:00:24.04" />
                    <SPLIT distance="75" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:00:51.23" />
                    <SPLIT distance="125" swimtime="00:01:05.18" />
                    <SPLIT distance="150" swimtime="00:01:19.76" />
                    <SPLIT distance="175" swimtime="00:01:35.10" />
                    <SPLIT distance="200" swimtime="00:01:50.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="21" place="1" lane="5" heat="3" heatid="30021" swimtime="00:01:49.93" reactiontime="+63" points="954">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.12" />
                    <SPLIT distance="50" swimtime="00:00:24.31" />
                    <SPLIT distance="75" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:00:51.69" />
                    <SPLIT distance="125" swimtime="00:01:05.93" />
                    <SPLIT distance="150" swimtime="00:01:20.43" />
                    <SPLIT distance="175" swimtime="00:01:34.93" />
                    <SPLIT distance="200" swimtime="00:01:49.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150418" lastname="SMITH" firstname="Kieran" gender="M" birthdate="2000-05-20">
              <ENTRIES>
                <ENTRY entrytime="00:01:41.78" eventid="44" heat="4" lane="5">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:03:35.99" eventid="24" heat="5" lane="4">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
                <ENTRY entrytime="NT" eventid="35" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="44" place="9" lane="5" heat="4" heatid="40044" swimtime="00:01:42.54" reactiontime="+68" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.13" />
                    <SPLIT distance="50" swimtime="00:00:23.87" />
                    <SPLIT distance="75" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:00:49.98" />
                    <SPLIT distance="125" swimtime="00:01:03.17" />
                    <SPLIT distance="150" swimtime="00:01:16.48" />
                    <SPLIT distance="175" swimtime="00:01:29.71" />
                    <SPLIT distance="200" swimtime="00:01:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="124" place="1" lane="4" heat="1" heatid="10124" swimtime="00:03:34.38" reactiontime="+68" points="970">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.33" />
                    <SPLIT distance="50" swimtime="00:00:24.41" />
                    <SPLIT distance="75" swimtime="00:00:37.68" />
                    <SPLIT distance="100" swimtime="00:00:51.07" />
                    <SPLIT distance="125" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:17.88" />
                    <SPLIT distance="175" swimtime="00:01:31.35" />
                    <SPLIT distance="200" swimtime="00:01:44.91" />
                    <SPLIT distance="225" swimtime="00:01:58.66" />
                    <SPLIT distance="250" swimtime="00:02:12.33" />
                    <SPLIT distance="275" swimtime="00:02:25.90" />
                    <SPLIT distance="300" swimtime="00:02:39.61" />
                    <SPLIT distance="325" swimtime="00:02:53.35" />
                    <SPLIT distance="350" swimtime="00:03:07.22" />
                    <SPLIT distance="375" swimtime="00:03:21.25" />
                    <SPLIT distance="400" swimtime="00:03:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="1" lane="4" heat="5" heatid="50024" swimtime="00:03:36.91" reactiontime="+69" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:24.91" />
                    <SPLIT distance="75" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:00:52.13" />
                    <SPLIT distance="125" swimtime="00:01:05.81" />
                    <SPLIT distance="150" swimtime="00:01:19.48" />
                    <SPLIT distance="175" swimtime="00:01:33.20" />
                    <SPLIT distance="200" swimtime="00:01:46.96" />
                    <SPLIT distance="225" swimtime="00:02:00.79" />
                    <SPLIT distance="250" swimtime="00:02:14.48" />
                    <SPLIT distance="275" swimtime="00:02:28.33" />
                    <SPLIT distance="300" swimtime="00:02:42.08" />
                    <SPLIT distance="325" swimtime="00:02:56.01" />
                    <SPLIT distance="350" swimtime="00:03:09.86" />
                    <SPLIT distance="375" swimtime="00:03:23.77" />
                    <SPLIT distance="400" swimtime="00:03:36.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150412" lastname="FOSTER" firstname="Carson" gender="M" birthdate="2001-10-26">
              <ENTRIES>
                <ENTRY entrytime="00:01:51.35" eventid="7" heat="5" lane="5">
                  <MEETINFO date="2021-12-16" />
                </ENTRY>
                <ENTRY entrytime="00:03:57.99" eventid="37" heat="2" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="48" />
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="107" place="2" lane="5" heat="1" heatid="10107" swimtime="00:01:50.96" reactiontime="+67" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.02" />
                    <SPLIT distance="50" swimtime="00:00:24.10" />
                    <SPLIT distance="75" swimtime="00:00:38.08" />
                    <SPLIT distance="100" swimtime="00:00:51.36" />
                    <SPLIT distance="125" swimtime="00:01:07.59" />
                    <SPLIT distance="150" swimtime="00:01:24.06" />
                    <SPLIT distance="175" swimtime="00:01:38.12" />
                    <SPLIT distance="200" swimtime="00:01:50.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="2" lane="5" heat="5" heatid="50007" swimtime="00:01:51.89" reactiontime="+66" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.99" />
                    <SPLIT distance="50" swimtime="00:00:24.04" />
                    <SPLIT distance="75" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:00:51.60" />
                    <SPLIT distance="125" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:24.11" />
                    <SPLIT distance="175" swimtime="00:01:38.68" />
                    <SPLIT distance="200" swimtime="00:01:51.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="137" place="2" lane="5" heat="1" heatid="10137" swimtime="00:03:57.63" reactiontime="+69" points="964">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:25.10" />
                    <SPLIT distance="75" swimtime="00:00:39.45" />
                    <SPLIT distance="100" swimtime="00:00:53.92" />
                    <SPLIT distance="125" swimtime="00:01:09.22" />
                    <SPLIT distance="150" swimtime="00:01:23.80" />
                    <SPLIT distance="175" swimtime="00:01:38.49" />
                    <SPLIT distance="200" swimtime="00:01:53.01" />
                    <SPLIT distance="225" swimtime="00:02:09.77" />
                    <SPLIT distance="250" swimtime="00:02:26.91" />
                    <SPLIT distance="275" swimtime="00:02:44.10" />
                    <SPLIT distance="300" swimtime="00:03:01.30" />
                    <SPLIT distance="325" swimtime="00:03:15.97" />
                    <SPLIT distance="350" swimtime="00:03:29.68" />
                    <SPLIT distance="375" swimtime="00:03:43.81" />
                    <SPLIT distance="400" swimtime="00:03:57.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="2" lane="4" heat="2" heatid="20037" swimtime="00:04:01.34" reactiontime="+67" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.67" />
                    <SPLIT distance="50" swimtime="00:00:25.67" />
                    <SPLIT distance="75" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:00:54.68" />
                    <SPLIT distance="125" swimtime="00:01:10.03" />
                    <SPLIT distance="150" swimtime="00:01:24.74" />
                    <SPLIT distance="175" swimtime="00:01:39.54" />
                    <SPLIT distance="200" swimtime="00:01:53.98" />
                    <SPLIT distance="225" swimtime="00:02:11.01" />
                    <SPLIT distance="250" swimtime="00:02:28.05" />
                    <SPLIT distance="275" swimtime="00:02:45.22" />
                    <SPLIT distance="300" swimtime="00:03:02.34" />
                    <SPLIT distance="325" swimtime="00:03:17.76" />
                    <SPLIT distance="350" swimtime="00:03:32.18" />
                    <SPLIT distance="375" swimtime="00:03:47.05" />
                    <SPLIT distance="400" swimtime="00:04:01.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183501" lastname="MAGAHEY" firstname="Jake" gender="M" birthdate="2001-09-14">
              <ENTRIES>
                <ENTRY entrytime="00:03:38.02" eventid="24" heat="5" lane="6">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="124" place="7" lane="8" heat="1" heatid="10124" swimtime="00:03:38.12" reactiontime="+74" points="921">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.76" />
                    <SPLIT distance="50" swimtime="00:00:25.26" />
                    <SPLIT distance="75" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:00:52.91" />
                    <SPLIT distance="125" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:20.61" />
                    <SPLIT distance="175" swimtime="00:01:34.44" />
                    <SPLIT distance="200" swimtime="00:01:48.51" />
                    <SPLIT distance="225" swimtime="00:02:02.29" />
                    <SPLIT distance="250" swimtime="00:02:16.26" />
                    <SPLIT distance="275" swimtime="00:02:30.00" />
                    <SPLIT distance="300" swimtime="00:02:43.95" />
                    <SPLIT distance="325" swimtime="00:02:57.51" />
                    <SPLIT distance="350" swimtime="00:03:11.43" />
                    <SPLIT distance="375" swimtime="00:03:25.05" />
                    <SPLIT distance="400" swimtime="00:03:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="24" place="8" lane="6" heat="5" heatid="50024" swimtime="00:03:38.74" reactiontime="+74" points="913">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.11" />
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                    <SPLIT distance="75" swimtime="00:00:39.49" />
                    <SPLIT distance="100" swimtime="00:00:53.47" />
                    <SPLIT distance="125" swimtime="00:01:07.30" />
                    <SPLIT distance="150" swimtime="00:01:21.19" />
                    <SPLIT distance="175" swimtime="00:01:35.05" />
                    <SPLIT distance="200" swimtime="00:01:49.00" />
                    <SPLIT distance="225" swimtime="00:02:02.88" />
                    <SPLIT distance="250" swimtime="00:02:16.66" />
                    <SPLIT distance="275" swimtime="00:02:30.27" />
                    <SPLIT distance="300" swimtime="00:02:43.98" />
                    <SPLIT distance="325" swimtime="00:02:57.46" />
                    <SPLIT distance="350" swimtime="00:03:11.30" />
                    <SPLIT distance="375" swimtime="00:03:25.12" />
                    <SPLIT distance="400" swimtime="00:03:38.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="214519" lastname="FOSTER" firstname="Jake" gender="M" birthdate="2000-09-06">
              <ENTRIES>
                <ENTRY entrytime="00:04:13.76" eventid="37" heat="1" lane="4">
                  <MEETINFO date="2022-04-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="32" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="137" place="6" lane="6" heat="1" heatid="10137" swimtime="00:04:02.51" reactiontime="+65" points="907">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.58" />
                    <SPLIT distance="50" swimtime="00:00:25.44" />
                    <SPLIT distance="75" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:00:54.95" />
                    <SPLIT distance="125" swimtime="00:01:11.04" />
                    <SPLIT distance="150" swimtime="00:01:26.55" />
                    <SPLIT distance="175" swimtime="00:01:42.29" />
                    <SPLIT distance="200" swimtime="00:01:57.84" />
                    <SPLIT distance="225" swimtime="00:02:14.20" />
                    <SPLIT distance="250" swimtime="00:02:30.94" />
                    <SPLIT distance="275" swimtime="00:02:47.89" />
                    <SPLIT distance="300" swimtime="00:03:05.14" />
                    <SPLIT distance="325" swimtime="00:03:20.27" />
                    <SPLIT distance="350" swimtime="00:03:34.80" />
                    <SPLIT distance="375" swimtime="00:03:49.02" />
                    <SPLIT distance="400" swimtime="00:04:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="37" place="4" lane="4" heat="1" heatid="10037" swimtime="00:04:02.64" reactiontime="+64" points="906">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.85" />
                    <SPLIT distance="50" swimtime="00:00:25.88" />
                    <SPLIT distance="75" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:00:55.35" />
                    <SPLIT distance="125" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:26.97" />
                    <SPLIT distance="175" swimtime="00:01:42.54" />
                    <SPLIT distance="200" swimtime="00:01:57.90" />
                    <SPLIT distance="225" swimtime="00:02:14.12" />
                    <SPLIT distance="250" swimtime="00:02:30.89" />
                    <SPLIT distance="275" swimtime="00:02:47.91" />
                    <SPLIT distance="300" swimtime="00:03:04.97" />
                    <SPLIT distance="325" swimtime="00:03:20.09" />
                    <SPLIT distance="350" swimtime="00:03:34.45" />
                    <SPLIT distance="375" swimtime="00:03:48.84" />
                    <SPLIT distance="400" swimtime="00:04:02.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183484" lastname="CURTISS" firstname="David" gender="M" birthdate="2002-07-04">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="9" />
                <ENTRY entrytime="NT" eventid="26" />
                <ENTRY entrytime="00:00:21.84" eventid="31" heat="7" lane="4">
                  <MEETINFO date="2022-08-21" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="27" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="31" place="24" lane="4" heat="7" heatid="70031" swimtime="00:00:21.40" reactiontime="+63" points="836">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.27" />
                    <SPLIT distance="50" swimtime="00:00:21.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183566" lastname="CURZAN" firstname="Claire" gender="F" birthdate="2004-06-30">
              <ENTRIES>
                <ENTRY entrytime="00:00:58.39" eventid="2" heat="5" lane="1">
                  <MEETINFO date="2022-04-29" />
                </ENTRY>
                <ENTRY entrytime="00:00:55.39" eventid="38" heat="2" lane="4">
                  <MEETINFO date="2021-12-21" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.31" eventid="45" heat="3" lane="1">
                  <MEETINFO date="2022-03-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:28.09" eventid="18" heat="4" lane="5">
                  <MEETINFO date="2022-04-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.55" eventid="4" heat="6" lane="4">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:23.80" eventid="30" heat="6" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="3" lane="3" heat="1" heatid="10102" swimtime="00:00:55.74" reactiontime="+59" points="954">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                    <SPLIT distance="75" swimtime="00:00:41.19" />
                    <SPLIT distance="100" swimtime="00:00:55.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="9" lane="1" heat="5" heatid="50002" swimtime="00:00:56.90" reactiontime="+60" points="897">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                    <SPLIT distance="50" swimtime="00:00:27.46" />
                    <SPLIT distance="75" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:00:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="3" lane="2" heat="2" heatid="20202" swimtime="00:00:56.08" reactiontime="+61" points="937">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.08" />
                    <SPLIT distance="50" swimtime="00:00:27.02" />
                    <SPLIT distance="75" swimtime="00:00:41.59" />
                    <SPLIT distance="100" swimtime="00:00:56.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="10" lane="4" heat="2" heatid="20038" swimtime="00:00:56.90" reactiontime="+55" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:26.05" />
                    <SPLIT distance="75" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:00:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="5" lane="2" heat="1" heatid="10238" swimtime="00:00:56.37" reactiontime="+64" points="908">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.93" />
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                    <SPLIT distance="75" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:00:56.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="145" place="2" lane="4" heat="1" heatid="10145" swimtime="00:02:00.53" reactiontime="+59" points="960">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="75" swimtime="00:00:43.39" />
                    <SPLIT distance="100" swimtime="00:00:58.39" />
                    <SPLIT distance="125" swimtime="00:01:13.84" />
                    <SPLIT distance="150" swimtime="00:01:29.25" />
                    <SPLIT distance="175" swimtime="00:01:44.91" />
                    <SPLIT distance="200" swimtime="00:02:00.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="1" lane="1" heat="3" heatid="30045" swimtime="00:02:02.05" reactiontime="+60" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.50" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                    <SPLIT distance="75" swimtime="00:00:43.49" />
                    <SPLIT distance="100" swimtime="00:00:58.96" />
                    <SPLIT distance="125" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:30.08" />
                    <SPLIT distance="175" swimtime="00:01:46.13" />
                    <SPLIT distance="200" swimtime="00:02:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="118" place="2" lane="4" heat="1" heatid="10118" swimtime="00:00:25.54" reactiontime="+60" points="968">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.54" />
                    <SPLIT distance="50" swimtime="00:00:25.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="4" lane="5" heat="4" heatid="40018" swimtime="00:00:26.07" reactiontime="+60" points="910">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.75" />
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="1" lane="5" heat="1" heatid="10218" swimtime="00:00:25.60" reactiontime="+60" points="961">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.61" />
                    <SPLIT distance="50" swimtime="00:00:25.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="104" place="5" lane="7" heat="1" heatid="10104" swimtime="00:00:24.92" reactiontime="+62" points="936">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.41" />
                    <SPLIT distance="50" swimtime="00:00:24.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="11" lane="4" heat="6" heatid="60004" swimtime="00:00:25.43" reactiontime="+67" points="881">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="6" lane="7" heat="2" heatid="20204" swimtime="00:00:24.96" reactiontime="+64" points="931">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:24.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="10" lane="4" heat="6" heatid="60030" swimtime="00:00:24.17" reactiontime="+60" points="853">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.66" />
                    <SPLIT distance="50" swimtime="00:00:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="12" lane="2" heat="1" heatid="10230" swimtime="00:00:24.22" reactiontime="+60" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.61" />
                    <SPLIT distance="50" swimtime="00:00:24.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="197516" lastname="STADDEN" firstname="Isabelle" gender="F" birthdate="2002-07-09">
              <ENTRIES>
                <ENTRY entrytime="00:00:59.16" eventid="2" heat="4" lane="8">
                  <MEETINFO date="2022-04-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:02.20" eventid="45" heat="3" lane="5">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="102" place="8" lane="1" heat="1" heatid="10102" swimtime="00:00:57.20" reactiontime="+60" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.44" />
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                    <SPLIT distance="75" swimtime="00:00:42.29" />
                    <SPLIT distance="100" swimtime="00:00:57.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2" place="7" lane="8" heat="4" heatid="40002" swimtime="00:00:56.85" reactiontime="+61" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.45" />
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="75" swimtime="00:00:42.33" />
                    <SPLIT distance="100" swimtime="00:00:56.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="202" place="7" lane="6" heat="2" heatid="20202" swimtime="00:00:56.45" reactiontime="+59" points="919">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.39" />
                    <SPLIT distance="50" swimtime="00:00:27.39" />
                    <SPLIT distance="75" swimtime="00:00:42.04" />
                    <SPLIT distance="100" swimtime="00:00:56.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="45" place="9" lane="5" heat="3" heatid="30045" swimtime="00:02:03.78" reactiontime="+66" points="887">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.96" />
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="75" swimtime="00:00:44.45" />
                    <SPLIT distance="100" swimtime="00:01:00.11" />
                    <SPLIT distance="125" swimtime="00:01:16.51" />
                    <SPLIT distance="150" swimtime="00:01:32.34" />
                    <SPLIT distance="175" swimtime="00:01:48.22" />
                    <SPLIT distance="200" swimtime="00:02:03.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="130153" lastname="KING" firstname="Lilly" gender="F" birthdate="1997-02-10">
              <ENTRIES>
                <ENTRY entrytime="00:01:03.23" eventid="15" heat="5" lane="4">
                  <MEETINFO date="2022-10-29" />
                </ENTRY>
                <ENTRY entrytime="00:02:16.47" eventid="28" heat="5" lane="4">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="00:00:29.15" eventid="40" heat="6" lane="4">
                  <MEETINFO date="2021-09-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="115" place="1" lane="4" heat="1" heatid="10115" swimtime="00:01:02.67" reactiontime="+63" points="985">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.48" />
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="75" swimtime="00:00:45.77" />
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="15" place="3" lane="4" heat="5" heatid="50015" swimtime="00:01:03.94" reactiontime="+63" points="927">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="75" swimtime="00:00:46.81" />
                    <SPLIT distance="100" swimtime="00:01:03.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="215" place="1" lane="5" heat="2" heatid="20215" swimtime="00:01:03.33" reactiontime="+64" points="954">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                    <SPLIT distance="75" swimtime="00:00:46.45" />
                    <SPLIT distance="100" swimtime="00:01:03.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="128" place="2" lane="5" heat="1" heatid="10128" swimtime="00:02:17.13" reactiontime="+64" points="945">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.73" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:47.71" />
                    <SPLIT distance="100" swimtime="00:01:05.23" />
                    <SPLIT distance="125" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:01:41.00" />
                    <SPLIT distance="175" swimtime="00:01:59.04" />
                    <SPLIT distance="200" swimtime="00:02:17.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="2" lane="4" heat="5" heatid="50028" swimtime="00:02:18.59" reactiontime="+65" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.79" />
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="75" swimtime="00:00:48.31" />
                    <SPLIT distance="100" swimtime="00:01:06.12" />
                    <SPLIT distance="125" swimtime="00:01:24.52" />
                    <SPLIT distance="150" swimtime="00:01:43.42" />
                    <SPLIT distance="175" swimtime="00:02:01.13" />
                    <SPLIT distance="200" swimtime="00:02:18.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="140" place="3" lane="5" heat="1" heatid="10140" swimtime="00:00:29.11" reactiontime="+62" points="944">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.33" />
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="5" lane="4" heat="6" heatid="60040" swimtime="00:00:29.53" reactiontime="+62" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="240" place="2" lane="3" heat="2" heatid="20240" swimtime="00:00:28.86" reactiontime="+64" points="969">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.30" />
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="156655" lastname="LAZOR" firstname="Annie" gender="F" birthdate="1994-08-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:04.83" eventid="15" heat="6" lane="6">
                  <MEETINFO date="2021-11-14" />
                </ENTRY>
                <ENTRY entrytime="00:00:30.89" eventid="40" heat="4" lane="3">
                  <MEETINFO date="2022-06-24" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="15" place="20" lane="6" heat="6" heatid="60015" swimtime="00:01:05.51" reactiontime="+71" points="862">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="75" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="40" place="23" lane="3" heat="4" heatid="40040" swimtime="00:00:30.69" reactiontime="+68" points="805">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.18" />
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183578" lastname="HUSKE" firstname="Torri" gender="F" birthdate="2002-12-07">
              <ENTRIES>
                <ENTRY entrytime="00:00:55.64" eventid="38" heat="3" lane="5">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="00:00:51.93" eventid="13" heat="8" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:24.88" eventid="4" heat="4" lane="4">
                  <MEETINFO date="2021-12-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="138" place="2" lane="4" heat="1" heatid="10138" swimtime="00:00:54.75" reactiontime="+59" points="991">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.48" />
                    <SPLIT distance="50" swimtime="00:00:25.08" />
                    <SPLIT distance="75" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:00:54.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="38" place="2" lane="5" heat="3" heatid="30038" swimtime="00:00:56.01" reactiontime="+59" points="925">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.62" />
                    <SPLIT distance="50" swimtime="00:00:25.50" />
                    <SPLIT distance="75" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="238" place="1" lane="4" heat="1" heatid="10238" swimtime="00:00:55.23" reactiontime="+60" points="965">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.56" />
                    <SPLIT distance="50" swimtime="00:00:25.48" />
                    <SPLIT distance="75" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:00:55.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="113" place="5" lane="7" heat="1" heatid="10113" swimtime="00:00:52.04" reactiontime="+62" points="900">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.59" />
                    <SPLIT distance="50" swimtime="00:00:24.68" />
                    <SPLIT distance="75" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:00:52.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="6" lane="3" heat="8" heatid="80013" swimtime="00:00:52.48" reactiontime="+63" points="877">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.69" />
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="75" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="6" lane="3" heat="1" heatid="10213" swimtime="00:00:52.11" reactiontime="+61" points="896">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.70" />
                    <SPLIT distance="50" swimtime="00:00:24.80" />
                    <SPLIT distance="75" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="104" place="1" lane="3" heat="1" heatid="10104" swimtime="00:00:24.64" reactiontime="+59" points="968">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.26" />
                    <SPLIT distance="50" swimtime="00:00:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4" place="4" lane="4" heat="4" heatid="40004" swimtime="00:00:25.11" reactiontime="+63" points="915">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.47" />
                    <SPLIT distance="50" swimtime="00:00:25.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="204" place="3" lane="5" heat="1" heatid="10204" swimtime="00:00:24.86" reactiontime="+61" points="943">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.27" />
                    <SPLIT distance="50" swimtime="00:00:24.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="202573" lastname="HINDS" firstname="Natalie" gender="F" birthdate="1993-12-07">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:00:52.02" eventid="13" heat="8" lane="6">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="113" place="8" lane="1" heat="1" heatid="10113" swimtime="00:00:52.24" reactiontime="+65" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:24.90" />
                    <SPLIT distance="75" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:00:52.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="13" place="11" lane="6" heat="8" heatid="80013" swimtime="00:00:52.86" reactiontime="+67" points="859">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.97" />
                    <SPLIT distance="50" swimtime="00:00:25.24" />
                    <SPLIT distance="75" swimtime="00:00:38.95" />
                    <SPLIT distance="100" swimtime="00:00:52.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="213" place="7" lane="7" heat="2" heatid="20213" swimtime="00:00:52.16" reactiontime="+67" points="894">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.75" />
                    <SPLIT distance="50" swimtime="00:00:24.88" />
                    <SPLIT distance="75" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:00:52.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150313" lastname="DOUGLASS" firstname="Kate" gender="F" birthdate="2001-11-17">
              <ENTRIES>
                <ENTRY entrytime="00:02:21.43" eventid="28" heat="4" lane="7">
                  <MEETINFO date="2022-04-27" />
                </ENTRY>
                <ENTRY entrytime="00:02:04.24" eventid="6" heat="5" lane="4">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="128" place="1" lane="4" heat="1" heatid="10128" swimtime="00:02:15.77" reactiontime="+65" points="973">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                    <SPLIT distance="75" swimtime="00:00:48.02" />
                    <SPLIT distance="100" swimtime="00:01:05.35" />
                    <SPLIT distance="125" swimtime="00:01:23.01" />
                    <SPLIT distance="150" swimtime="00:01:40.65" />
                    <SPLIT distance="175" swimtime="00:01:58.19" />
                    <SPLIT distance="200" swimtime="00:02:15.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="28" place="1" lane="7" heat="4" heatid="40028" swimtime="00:02:16.52" reactiontime="+67" points="957">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="75" swimtime="00:00:48.48" />
                    <SPLIT distance="100" swimtime="00:01:05.82" />
                    <SPLIT distance="125" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:01:41.09" />
                    <SPLIT distance="175" swimtime="00:01:58.79" />
                    <SPLIT distance="200" swimtime="00:02:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="106" place="1" lane="4" heat="1" heatid="10106" swimtime="00:02:02.12" reactiontime="+67" points="993">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.99" />
                    <SPLIT distance="50" swimtime="00:00:26.34" />
                    <SPLIT distance="75" swimtime="00:00:42.35" />
                    <SPLIT distance="100" swimtime="00:00:57.63" />
                    <SPLIT distance="125" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:01:32.99" />
                    <SPLIT distance="175" swimtime="00:01:48.15" />
                    <SPLIT distance="200" swimtime="00:02:02.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="1" lane="4" heat="5" heatid="50006" swimtime="00:02:04.39" reactiontime="+67" points="940">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.02" />
                    <SPLIT distance="50" swimtime="00:00:26.49" />
                    <SPLIT distance="75" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:00:58.32" />
                    <SPLIT distance="125" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:33.97" />
                    <SPLIT distance="175" swimtime="00:01:49.85" />
                    <SPLIT distance="200" swimtime="00:02:04.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124875" lastname="LUTHER" firstname="Dakota" gender="F" birthdate="1999-11-07">
              <ENTRIES>
                <ENTRY entrytime="00:02:07.02" eventid="20" heat="4" lane="2">
                  <MEETINFO date="2022-07-26" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="120" place="1" lane="4" heat="1" heatid="10120" swimtime="00:02:03.37" reactiontime="+74" points="911">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="75" swimtime="00:00:43.23" />
                    <SPLIT distance="100" swimtime="00:00:58.94" />
                    <SPLIT distance="125" swimtime="00:01:14.85" />
                    <SPLIT distance="150" swimtime="00:01:30.97" />
                    <SPLIT distance="175" swimtime="00:01:47.13" />
                    <SPLIT distance="200" swimtime="00:02:03.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="1" lane="2" heat="4" heatid="40020" swimtime="00:02:03.73" reactiontime="+71" points="903">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.82" />
                    <SPLIT distance="50" swimtime="00:00:27.83" />
                    <SPLIT distance="75" swimtime="00:00:43.42" />
                    <SPLIT distance="100" swimtime="00:00:59.16" />
                    <SPLIT distance="125" swimtime="00:01:14.95" />
                    <SPLIT distance="150" swimtime="00:01:31.00" />
                    <SPLIT distance="175" swimtime="00:01:47.31" />
                    <SPLIT distance="200" swimtime="00:02:03.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="143364" lastname="FLICKINGER" firstname="Hali" gender="F" birthdate="1994-07-07">
              <ENTRIES>
                <ENTRY entrytime="00:02:03.73" eventid="20" heat="3" lane="4">
                  <MEETINFO date="2021-12-04" />
                </ENTRY>
                <ENTRY entrytime="00:01:54.36" eventid="43" heat="5" lane="6">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
                <ENTRY entrytime="00:04:29.82" eventid="36" heat="4" lane="3">
                  <MEETINFO date="2021-11-28" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="120" place="2" lane="5" heat="1" heatid="10120" swimtime="00:02:03.78" reactiontime="+69" points="902">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="75" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:00:58.82" />
                    <SPLIT distance="125" swimtime="00:01:14.66" />
                    <SPLIT distance="150" swimtime="00:01:30.84" />
                    <SPLIT distance="175" swimtime="00:01:47.32" />
                    <SPLIT distance="200" swimtime="00:02:03.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="20" place="2" lane="4" heat="3" heatid="30020" swimtime="00:02:04.66" reactiontime="+71" points="883">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.17" />
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="75" swimtime="00:00:44.17" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="125" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:01:31.99" />
                    <SPLIT distance="175" swimtime="00:01:48.31" />
                    <SPLIT distance="200" swimtime="00:02:04.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="9" lane="6" heat="5" heatid="50043" swimtime="00:01:54.20" reactiontime="+67" points="901">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="75" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:00:55.99" />
                    <SPLIT distance="125" swimtime="00:01:10.52" />
                    <SPLIT distance="150" swimtime="00:01:25.30" />
                    <SPLIT distance="175" swimtime="00:01:39.94" />
                    <SPLIT distance="200" swimtime="00:01:54.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="1" lane="2" heat="1" heatid="10136" swimtime="00:04:26.51" reactiontime="+59" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:44.07" />
                    <SPLIT distance="100" swimtime="00:01:00.06" />
                    <SPLIT distance="125" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:01:34.10" />
                    <SPLIT distance="175" swimtime="00:01:50.48" />
                    <SPLIT distance="200" swimtime="00:02:06.97" />
                    <SPLIT distance="225" swimtime="00:02:26.61" />
                    <SPLIT distance="250" swimtime="00:02:46.27" />
                    <SPLIT distance="275" swimtime="00:03:05.99" />
                    <SPLIT distance="300" swimtime="00:03:25.72" />
                    <SPLIT distance="325" swimtime="00:03:41.55" />
                    <SPLIT distance="350" swimtime="00:03:56.62" />
                    <SPLIT distance="375" swimtime="00:04:11.76" />
                    <SPLIT distance="400" swimtime="00:04:26.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="5" lane="3" heat="4" heatid="40036" swimtime="00:04:31.61" reactiontime="+68" points="866">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="75" swimtime="00:00:44.57" />
                    <SPLIT distance="100" swimtime="00:01:00.75" />
                    <SPLIT distance="125" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:01:35.50" />
                    <SPLIT distance="175" swimtime="00:01:52.40" />
                    <SPLIT distance="200" swimtime="00:02:09.18" />
                    <SPLIT distance="225" swimtime="00:02:28.97" />
                    <SPLIT distance="250" swimtime="00:02:48.98" />
                    <SPLIT distance="275" swimtime="00:03:08.91" />
                    <SPLIT distance="300" swimtime="00:03:28.85" />
                    <SPLIT distance="325" swimtime="00:03:45.34" />
                    <SPLIT distance="350" swimtime="00:04:00.94" />
                    <SPLIT distance="375" swimtime="00:04:16.38" />
                    <SPLIT distance="400" swimtime="00:04:31.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="183572" lastname="GEMMELL" firstname="Erin" gender="F" birthdate="2004-12-02">
              <ENTRIES>
                <ENTRY entrytime="00:01:53.27" eventid="43" heat="4" lane="3">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="00:04:00.45" eventid="1" heat="4" lane="3">
                  <MEETINFO date="2022-11-03" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="143" place="4" lane="3" heat="1" heatid="10143" swimtime="00:01:52.56" reactiontime="+80" points="941">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.35" />
                    <SPLIT distance="75" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:00:55.18" />
                    <SPLIT distance="125" swimtime="00:01:09.48" />
                    <SPLIT distance="150" swimtime="00:01:24.11" />
                    <SPLIT distance="175" swimtime="00:01:38.51" />
                    <SPLIT distance="200" swimtime="00:01:52.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="43" place="3" lane="3" heat="4" heatid="40043" swimtime="00:01:53.47" reactiontime="+78" points="918">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                    <SPLIT distance="75" swimtime="00:00:40.91" />
                    <SPLIT distance="100" swimtime="00:00:55.44" />
                    <SPLIT distance="125" swimtime="00:01:09.94" />
                    <SPLIT distance="150" swimtime="00:01:24.62" />
                    <SPLIT distance="175" swimtime="00:01:39.21" />
                    <SPLIT distance="200" swimtime="00:01:53.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="101" place="6" lane="3" heat="1" heatid="10101" swimtime="00:04:01.82" reactiontime="+80" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.12" />
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                    <SPLIT distance="75" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:00:57.13" />
                    <SPLIT distance="125" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:27.62" />
                    <SPLIT distance="175" swimtime="00:01:43.00" />
                    <SPLIT distance="200" swimtime="00:01:58.48" />
                    <SPLIT distance="225" swimtime="00:02:13.94" />
                    <SPLIT distance="250" swimtime="00:02:29.58" />
                    <SPLIT distance="275" swimtime="00:02:45.42" />
                    <SPLIT distance="300" swimtime="00:03:01.27" />
                    <SPLIT distance="325" swimtime="00:03:16.77" />
                    <SPLIT distance="350" swimtime="00:03:32.27" />
                    <SPLIT distance="375" swimtime="00:03:47.25" />
                    <SPLIT distance="400" swimtime="00:04:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="3" lane="3" heat="4" heatid="40001" swimtime="00:04:00.49" reactiontime="+82" points="920">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.76" />
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="75" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:00:56.71" />
                    <SPLIT distance="125" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:27.03" />
                    <SPLIT distance="175" swimtime="00:01:42.26" />
                    <SPLIT distance="200" swimtime="00:01:57.63" />
                    <SPLIT distance="225" swimtime="00:02:12.82" />
                    <SPLIT distance="250" swimtime="00:02:28.10" />
                    <SPLIT distance="275" swimtime="00:02:43.40" />
                    <SPLIT distance="300" swimtime="00:02:58.96" />
                    <SPLIT distance="325" swimtime="00:03:14.41" />
                    <SPLIT distance="350" swimtime="00:03:30.22" />
                    <SPLIT distance="375" swimtime="00:03:45.43" />
                    <SPLIT distance="400" swimtime="00:04:00.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="150328" lastname="WALSH" firstname="Alex" gender="F" birthdate="2001-07-31">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="00:02:07.13" eventid="6" heat="3" lane="3">
                  <MEETINFO date="2022-06-19" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="NT" eventid="34" />
                <ENTRY entrytime="NT" eventid="11" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="106" place="2" lane="5" heat="1" heatid="10106" swimtime="00:02:03.37" reactiontime="+75" points="963">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.22" />
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                    <SPLIT distance="75" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:00:57.38" />
                    <SPLIT distance="125" swimtime="00:01:15.00" />
                    <SPLIT distance="150" swimtime="00:01:33.17" />
                    <SPLIT distance="175" swimtime="00:01:48.79" />
                    <SPLIT distance="200" swimtime="00:02:03.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6" place="2" lane="3" heat="3" heatid="30006" swimtime="00:02:05.94" reactiontime="+75" points="905">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                    <SPLIT distance="75" swimtime="00:00:43.57" />
                    <SPLIT distance="100" swimtime="00:00:58.72" />
                    <SPLIT distance="125" swimtime="00:01:16.76" />
                    <SPLIT distance="150" swimtime="00:01:35.03" />
                    <SPLIT distance="175" swimtime="00:01:51.45" />
                    <SPLIT distance="200" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="105648" lastname="SMITH" firstname="Leah" gender="F" birthdate="1995-04-19">
              <ENTRIES>
                <ENTRY entrytime="00:04:02.08" eventid="1" heat="3" lane="6">
                  <MEETINFO date="2022-06-18" />
                </ENTRY>
                <ENTRY entrytime="00:04:33.24" eventid="36" heat="4" lane="7">
                  <MEETINFO date="2022-11-04" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:08:12.01" eventid="12" heat="0" lane="2147483647">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="101" place="3" lane="6" heat="1" heatid="10101" swimtime="00:03:59.78" reactiontime="+71" points="928">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                    <SPLIT distance="75" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:00:57.82" />
                    <SPLIT distance="125" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:01:28.05" />
                    <SPLIT distance="175" swimtime="00:01:43.19" />
                    <SPLIT distance="200" swimtime="00:01:58.49" />
                    <SPLIT distance="225" swimtime="00:02:13.71" />
                    <SPLIT distance="250" swimtime="00:02:29.09" />
                    <SPLIT distance="275" swimtime="00:02:44.26" />
                    <SPLIT distance="300" swimtime="00:02:59.60" />
                    <SPLIT distance="325" swimtime="00:03:14.63" />
                    <SPLIT distance="350" swimtime="00:03:29.94" />
                    <SPLIT distance="375" swimtime="00:03:45.08" />
                    <SPLIT distance="400" swimtime="00:03:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1" place="4" lane="6" heat="3" heatid="30001" swimtime="00:04:00.71" reactiontime="+72" points="917">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:28.27" />
                    <SPLIT distance="75" swimtime="00:00:43.16" />
                    <SPLIT distance="100" swimtime="00:00:58.40" />
                    <SPLIT distance="125" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:28.94" />
                    <SPLIT distance="175" swimtime="00:01:44.04" />
                    <SPLIT distance="200" swimtime="00:01:59.40" />
                    <SPLIT distance="225" swimtime="00:02:14.60" />
                    <SPLIT distance="250" swimtime="00:02:30.00" />
                    <SPLIT distance="275" swimtime="00:02:45.18" />
                    <SPLIT distance="300" swimtime="00:03:00.44" />
                    <SPLIT distance="325" swimtime="00:03:15.49" />
                    <SPLIT distance="350" swimtime="00:03:30.86" />
                    <SPLIT distance="375" swimtime="00:03:46.14" />
                    <SPLIT distance="400" swimtime="00:04:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="136" place="4" lane="4" heat="1" heatid="10136" swimtime="00:04:29.18" reactiontime="+71" points="890">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.49" />
                    <SPLIT distance="50" swimtime="00:00:29.40" />
                    <SPLIT distance="75" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:02.96" />
                    <SPLIT distance="125" swimtime="00:01:20.83" />
                    <SPLIT distance="150" swimtime="00:01:37.54" />
                    <SPLIT distance="175" swimtime="00:01:54.40" />
                    <SPLIT distance="200" swimtime="00:02:11.06" />
                    <SPLIT distance="225" swimtime="00:02:30.18" />
                    <SPLIT distance="250" swimtime="00:02:49.65" />
                    <SPLIT distance="275" swimtime="00:03:09.41" />
                    <SPLIT distance="300" swimtime="00:03:29.36" />
                    <SPLIT distance="325" swimtime="00:03:45.13" />
                    <SPLIT distance="350" swimtime="00:03:59.96" />
                    <SPLIT distance="375" swimtime="00:04:14.86" />
                    <SPLIT distance="400" swimtime="00:04:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="36" place="1" lane="7" heat="4" heatid="40036" swimtime="00:04:30.93" reactiontime="+73" points="873">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.50" />
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="75" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:03.33" />
                    <SPLIT distance="125" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:01:37.92" />
                    <SPLIT distance="175" swimtime="00:01:54.78" />
                    <SPLIT distance="200" swimtime="00:02:11.57" />
                    <SPLIT distance="225" swimtime="00:02:30.78" />
                    <SPLIT distance="250" swimtime="00:02:50.32" />
                    <SPLIT distance="275" swimtime="00:03:10.08" />
                    <SPLIT distance="300" swimtime="00:03:30.00" />
                    <SPLIT distance="325" swimtime="00:03:46.10" />
                    <SPLIT distance="350" swimtime="00:04:01.32" />
                    <SPLIT distance="375" swimtime="00:04:16.38" />
                    <SPLIT distance="400" swimtime="00:04:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="112" place="4" lane="5" heat="5" heatid="30112" swimtime="00:08:14.24" reactiontime="+73" points="912">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.62" />
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                    <SPLIT distance="75" swimtime="00:00:43.70" />
                    <SPLIT distance="100" swimtime="00:00:59.09" />
                    <SPLIT distance="125" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:29.84" />
                    <SPLIT distance="175" swimtime="00:01:45.32" />
                    <SPLIT distance="200" swimtime="00:02:00.97" />
                    <SPLIT distance="225" swimtime="00:02:16.46" />
                    <SPLIT distance="250" swimtime="00:02:32.16" />
                    <SPLIT distance="275" swimtime="00:02:47.85" />
                    <SPLIT distance="300" swimtime="00:03:03.56" />
                    <SPLIT distance="325" swimtime="00:03:19.25" />
                    <SPLIT distance="350" swimtime="00:03:34.89" />
                    <SPLIT distance="375" swimtime="00:03:50.54" />
                    <SPLIT distance="400" swimtime="00:04:06.19" />
                    <SPLIT distance="425" swimtime="00:04:21.78" />
                    <SPLIT distance="450" swimtime="00:04:37.46" />
                    <SPLIT distance="475" swimtime="00:04:53.13" />
                    <SPLIT distance="500" swimtime="00:05:08.89" />
                    <SPLIT distance="525" swimtime="00:05:24.87" />
                    <SPLIT distance="550" swimtime="00:05:40.82" />
                    <SPLIT distance="575" swimtime="00:05:56.44" />
                    <SPLIT distance="600" swimtime="00:06:12.13" />
                    <SPLIT distance="625" swimtime="00:06:27.93" />
                    <SPLIT distance="650" swimtime="00:06:43.38" />
                    <SPLIT distance="675" swimtime="00:06:58.86" />
                    <SPLIT distance="700" swimtime="00:07:14.31" />
                    <SPLIT distance="725" swimtime="00:07:29.60" />
                    <SPLIT distance="750" swimtime="00:07:44.68" />
                    <SPLIT distance="775" swimtime="00:07:59.66" />
                    <SPLIT distance="800" swimtime="00:08:14.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="124845" lastname="BROWN" firstname="Erika" gender="F" birthdate="1998-08-27">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="27" />
                <ENTRY entrytime="NT" eventid="8" />
                <ENTRY entrytime="NT" eventid="47" />
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="NT" eventid="25" />
                <ENTRY entrytime="00:00:28.05" eventid="18" heat="4" lane="4">
                  <MEETINFO date="2022-04-28" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.02" eventid="30" heat="6" lane="6">
                  <MEETINFO date="2021-11-20" />
                </ENTRY>
                <ENTRY entrytime="NT" eventid="34" />
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="18" place="15" lane="4" heat="4" heatid="40018" swimtime="00:00:26.50" reactiontime="+60" points="867">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.16" />
                    <SPLIT distance="50" swimtime="00:00:26.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="218" place="16" lane="8" heat="2" heatid="20218" swimtime="00:00:26.56" reactiontime="+61" points="861">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.05" />
                    <SPLIT distance="50" swimtime="00:00:26.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="130" place="7" lane="1" heat="1" heatid="10130" swimtime="00:00:23.76" reactiontime="+59" points="898">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.52" />
                    <SPLIT distance="50" swimtime="00:00:23.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="8" lane="6" heat="6" heatid="60030" swimtime="00:00:23.98" reactiontime="+64" points="874">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.71" />
                    <SPLIT distance="50" swimtime="00:00:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="230" place="7" lane="6" heat="1" heatid="10230" swimtime="00:00:24.00" reactiontime="+65" points="872">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.65" />
                    <SPLIT distance="50" swimtime="00:00:24.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="213247" lastname="COX" firstname="Jillian" gender="F" birthdate="2005-07-18">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="17" />
                <ENTRY entrytime="00:08:22.94" eventid="12" heat="0" lane="-1">
                  <MEETINFO date="2022-11-05" />
                </ENTRY>
                <ENTRY entrytime="00:16:29.16" eventid="33" heat="2" lane="6">
                  <MEETINFO date="2022-08-27" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="112" place="6" lane="8" heat="5" heatid="30112" swimtime="00:08:20.95" reactiontime="+76" points="876">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.82" />
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                    <SPLIT distance="75" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:00:59.84" />
                    <SPLIT distance="125" swimtime="00:01:15.56" />
                    <SPLIT distance="150" swimtime="00:01:31.27" />
                    <SPLIT distance="175" swimtime="00:01:46.92" />
                    <SPLIT distance="200" swimtime="00:02:02.47" />
                    <SPLIT distance="225" swimtime="00:02:18.12" />
                    <SPLIT distance="250" swimtime="00:02:33.93" />
                    <SPLIT distance="275" swimtime="00:02:49.58" />
                    <SPLIT distance="300" swimtime="00:03:05.19" />
                    <SPLIT distance="325" swimtime="00:03:20.92" />
                    <SPLIT distance="350" swimtime="00:03:36.78" />
                    <SPLIT distance="375" swimtime="00:03:52.46" />
                    <SPLIT distance="400" swimtime="00:04:08.43" />
                    <SPLIT distance="425" swimtime="00:04:23.91" />
                    <SPLIT distance="450" swimtime="00:04:39.92" />
                    <SPLIT distance="475" swimtime="00:04:55.73" />
                    <SPLIT distance="500" swimtime="00:05:11.69" />
                    <SPLIT distance="525" swimtime="00:05:27.47" />
                    <SPLIT distance="550" swimtime="00:05:43.53" />
                    <SPLIT distance="575" swimtime="00:05:59.32" />
                    <SPLIT distance="600" swimtime="00:06:15.24" />
                    <SPLIT distance="625" swimtime="00:06:31.04" />
                    <SPLIT distance="650" swimtime="00:06:46.88" />
                    <SPLIT distance="675" swimtime="00:07:02.72" />
                    <SPLIT distance="700" swimtime="00:07:18.65" />
                    <SPLIT distance="725" swimtime="00:07:34.29" />
                    <SPLIT distance="750" swimtime="00:07:50.27" />
                    <SPLIT distance="775" swimtime="00:08:05.97" />
                    <SPLIT distance="800" swimtime="00:08:20.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="133" place="8" lane="6" heat="2" heatid="20033" swimtime="00:16:09.72" reactiontime="+67" points="848">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.52" />
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="75" swimtime="00:00:47.17" />
                    <SPLIT distance="100" swimtime="00:01:03.99" />
                    <SPLIT distance="125" swimtime="00:01:20.51" />
                    <SPLIT distance="150" swimtime="00:01:37.23" />
                    <SPLIT distance="175" swimtime="00:01:53.90" />
                    <SPLIT distance="200" swimtime="00:02:10.60" />
                    <SPLIT distance="225" swimtime="00:02:27.02" />
                    <SPLIT distance="250" swimtime="00:02:43.72" />
                    <SPLIT distance="275" swimtime="00:03:00.18" />
                    <SPLIT distance="300" swimtime="00:03:16.68" />
                    <SPLIT distance="325" swimtime="00:03:33.18" />
                    <SPLIT distance="350" swimtime="00:03:49.99" />
                    <SPLIT distance="375" swimtime="00:04:06.25" />
                    <SPLIT distance="400" swimtime="00:04:22.62" />
                    <SPLIT distance="425" swimtime="00:04:38.93" />
                    <SPLIT distance="450" swimtime="00:04:55.54" />
                    <SPLIT distance="475" swimtime="00:05:12.08" />
                    <SPLIT distance="500" swimtime="00:05:28.51" />
                    <SPLIT distance="525" swimtime="00:05:44.94" />
                    <SPLIT distance="550" swimtime="00:06:01.14" />
                    <SPLIT distance="575" swimtime="00:06:17.44" />
                    <SPLIT distance="600" swimtime="00:06:34.10" />
                    <SPLIT distance="625" swimtime="00:06:50.43" />
                    <SPLIT distance="650" swimtime="00:07:06.61" />
                    <SPLIT distance="675" swimtime="00:07:22.89" />
                    <SPLIT distance="700" swimtime="00:07:39.07" />
                    <SPLIT distance="725" swimtime="00:07:55.27" />
                    <SPLIT distance="750" swimtime="00:08:11.56" />
                    <SPLIT distance="775" swimtime="00:08:27.57" />
                    <SPLIT distance="800" swimtime="00:08:43.63" />
                    <SPLIT distance="825" swimtime="00:08:59.52" />
                    <SPLIT distance="850" swimtime="00:09:16.01" />
                    <SPLIT distance="875" swimtime="00:09:31.88" />
                    <SPLIT distance="900" swimtime="00:09:47.99" />
                    <SPLIT distance="925" swimtime="00:10:04.06" />
                    <SPLIT distance="950" swimtime="00:10:20.39" />
                    <SPLIT distance="975" swimtime="00:10:36.39" />
                    <SPLIT distance="1000" swimtime="00:10:52.48" />
                    <SPLIT distance="1025" swimtime="00:11:08.47" />
                    <SPLIT distance="1050" swimtime="00:11:24.56" />
                    <SPLIT distance="1075" swimtime="00:11:40.36" />
                    <SPLIT distance="1100" swimtime="00:11:56.55" />
                    <SPLIT distance="1125" swimtime="00:12:12.55" />
                    <SPLIT distance="1150" swimtime="00:12:28.80" />
                    <SPLIT distance="1175" swimtime="00:12:44.81" />
                    <SPLIT distance="1200" swimtime="00:13:00.86" />
                    <SPLIT distance="1225" swimtime="00:13:16.75" />
                    <SPLIT distance="1250" swimtime="00:13:32.65" />
                    <SPLIT distance="1275" swimtime="00:13:48.63" />
                    <SPLIT distance="1300" swimtime="00:14:04.74" />
                    <SPLIT distance="1325" swimtime="00:14:20.47" />
                    <SPLIT distance="1350" swimtime="00:14:36.49" />
                    <SPLIT distance="1375" swimtime="00:14:52.23" />
                    <SPLIT distance="1400" swimtime="00:15:08.15" />
                    <SPLIT distance="1425" swimtime="00:15:23.71" />
                    <SPLIT distance="1450" swimtime="00:15:39.46" />
                    <SPLIT distance="1475" swimtime="00:15:54.82" />
                    <SPLIT distance="1500" swimtime="00:16:09.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201580" lastname="MCMAHON" firstname="Kensey" gender="F" birthdate="1999-10-29">
              <ENTRIES>
                <ENTRY entrytime="00:16:16.22" eventid="33" heat="2" lane="5">
                  <MEETINFO date="2022-07-30" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="133" place="3" lane="5" heat="2" heatid="20033" swimtime="00:15:49.15" reactiontime="+75" points="904">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.59" />
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="75" swimtime="00:00:47.04" />
                    <SPLIT distance="100" swimtime="00:01:03.20" />
                    <SPLIT distance="125" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:01:35.40" />
                    <SPLIT distance="175" swimtime="00:01:51.44" />
                    <SPLIT distance="200" swimtime="00:02:07.51" />
                    <SPLIT distance="225" swimtime="00:02:23.40" />
                    <SPLIT distance="250" swimtime="00:02:39.20" />
                    <SPLIT distance="275" swimtime="00:02:55.13" />
                    <SPLIT distance="300" swimtime="00:03:10.93" />
                    <SPLIT distance="325" swimtime="00:03:26.61" />
                    <SPLIT distance="350" swimtime="00:03:42.29" />
                    <SPLIT distance="375" swimtime="00:03:58.11" />
                    <SPLIT distance="400" swimtime="00:04:13.81" />
                    <SPLIT distance="425" swimtime="00:04:29.66" />
                    <SPLIT distance="450" swimtime="00:04:45.39" />
                    <SPLIT distance="475" swimtime="00:05:01.18" />
                    <SPLIT distance="500" swimtime="00:05:16.85" />
                    <SPLIT distance="525" swimtime="00:05:32.45" />
                    <SPLIT distance="550" swimtime="00:05:48.01" />
                    <SPLIT distance="575" swimtime="00:06:03.65" />
                    <SPLIT distance="600" swimtime="00:06:19.28" />
                    <SPLIT distance="625" swimtime="00:06:34.94" />
                    <SPLIT distance="650" swimtime="00:06:50.62" />
                    <SPLIT distance="675" swimtime="00:07:06.36" />
                    <SPLIT distance="700" swimtime="00:07:22.13" />
                    <SPLIT distance="725" swimtime="00:07:37.92" />
                    <SPLIT distance="750" swimtime="00:07:53.75" />
                    <SPLIT distance="775" swimtime="00:08:09.51" />
                    <SPLIT distance="800" swimtime="00:08:25.42" />
                    <SPLIT distance="825" swimtime="00:08:41.40" />
                    <SPLIT distance="850" swimtime="00:08:57.38" />
                    <SPLIT distance="875" swimtime="00:09:13.34" />
                    <SPLIT distance="900" swimtime="00:09:29.13" />
                    <SPLIT distance="925" swimtime="00:09:44.98" />
                    <SPLIT distance="950" swimtime="00:10:00.91" />
                    <SPLIT distance="975" swimtime="00:10:16.64" />
                    <SPLIT distance="1000" swimtime="00:10:32.51" />
                    <SPLIT distance="1025" swimtime="00:10:48.31" />
                    <SPLIT distance="1050" swimtime="00:11:04.17" />
                    <SPLIT distance="1075" swimtime="00:11:20.02" />
                    <SPLIT distance="1100" swimtime="00:11:36.08" />
                    <SPLIT distance="1125" swimtime="00:11:52.05" />
                    <SPLIT distance="1150" swimtime="00:12:07.90" />
                    <SPLIT distance="1175" swimtime="00:12:23.91" />
                    <SPLIT distance="1200" swimtime="00:12:39.80" />
                    <SPLIT distance="1225" swimtime="00:12:55.62" />
                    <SPLIT distance="1250" swimtime="00:13:11.62" />
                    <SPLIT distance="1275" swimtime="00:13:27.69" />
                    <SPLIT distance="1300" swimtime="00:13:43.83" />
                    <SPLIT distance="1325" swimtime="00:13:59.51" />
                    <SPLIT distance="1350" swimtime="00:14:15.42" />
                    <SPLIT distance="1375" swimtime="00:14:31.20" />
                    <SPLIT distance="1400" swimtime="00:14:46.97" />
                    <SPLIT distance="1425" swimtime="00:15:02.87" />
                    <SPLIT distance="1450" swimtime="00:15:18.59" />
                    <SPLIT distance="1475" swimtime="00:15:34.26" />
                    <SPLIT distance="1500" swimtime="00:15:49.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="United States of America">
              <RESULTS>
                <RESULT eventid="109" place="3" lane="3" heat="1" swimtime="00:03:05.09" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.58" />
                    <SPLIT distance="50" swimtime="00:00:22.52" />
                    <SPLIT distance="75" swimtime="00:00:34.59" />
                    <SPLIT distance="100" swimtime="00:00:46.84" />
                    <SPLIT distance="125" swimtime="00:00:56.98" />
                    <SPLIT distance="150" swimtime="00:01:08.64" />
                    <SPLIT distance="175" swimtime="00:01:20.78" />
                    <SPLIT distance="200" swimtime="00:01:32.74" />
                    <SPLIT distance="225" swimtime="00:01:42.95" />
                    <SPLIT distance="250" swimtime="00:01:54.81" />
                    <SPLIT distance="275" swimtime="00:02:07.22" />
                    <SPLIT distance="300" swimtime="00:02:19.32" />
                    <SPLIT distance="325" swimtime="00:02:29.41" />
                    <SPLIT distance="350" swimtime="00:02:40.97" />
                    <SPLIT distance="375" swimtime="00:02:53.03" />
                    <SPLIT distance="400" swimtime="00:03:05.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="145806" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="197510" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="150412" reactiontime="+20" />
                    <RELAYPOSITION number="4" athleteid="150418" reactiontime="+27" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="9" place="3" lane="4" heat="1" swimtime="00:03:06.83" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.79" />
                    <SPLIT distance="50" swimtime="00:00:22.69" />
                    <SPLIT distance="75" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:00:48.07" />
                    <SPLIT distance="125" swimtime="00:00:58.11" />
                    <SPLIT distance="150" swimtime="00:01:09.82" />
                    <SPLIT distance="175" swimtime="00:01:21.81" />
                    <SPLIT distance="200" swimtime="00:01:33.98" />
                    <SPLIT distance="225" swimtime="00:01:44.31" />
                    <SPLIT distance="250" swimtime="00:01:55.94" />
                    <SPLIT distance="275" swimtime="00:02:08.27" />
                    <SPLIT distance="300" swimtime="00:02:20.75" />
                    <SPLIT distance="325" swimtime="00:02:30.81" />
                    <SPLIT distance="350" swimtime="00:02:42.61" />
                    <SPLIT distance="375" swimtime="00:02:54.77" />
                    <SPLIT distance="400" swimtime="00:03:06.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183484" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="145806" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="197514" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="150418" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="United States of America">
              <RESULTS>
                <RESULT eventid="148" place="1" lane="4" heat="1" swimtime="00:03:18.98" reactiontime="+54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.40" />
                    <SPLIT distance="50" swimtime="00:00:23.53" />
                    <SPLIT distance="75" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:00:48.96" />
                    <SPLIT distance="125" swimtime="00:01:00.17" />
                    <SPLIT distance="150" swimtime="00:01:14.13" />
                    <SPLIT distance="175" swimtime="00:01:28.78" />
                    <SPLIT distance="200" swimtime="00:01:43.84" />
                    <SPLIT distance="225" swimtime="00:01:53.87" />
                    <SPLIT distance="250" swimtime="00:02:06.40" />
                    <SPLIT distance="275" swimtime="00:02:19.48" />
                    <SPLIT distance="300" swimtime="00:02:33.03" />
                    <SPLIT distance="325" swimtime="00:02:43.12" />
                    <SPLIT distance="350" swimtime="00:02:54.81" />
                    <SPLIT distance="375" swimtime="00:03:06.94" />
                    <SPLIT distance="400" swimtime="00:03:18.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="105644" reactiontime="+54" />
                    <RELAYPOSITION number="2" athleteid="105614" reactiontime="+18" />
                    <RELAYPOSITION number="3" athleteid="197514" reactiontime="+15" />
                    <RELAYPOSITION number="4" athleteid="150418" reactiontime="+20" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="48" place="1" lane="4" heat="3" swimtime="00:03:23.55" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:24.35" />
                    <SPLIT distance="75" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:00:50.68" />
                    <SPLIT distance="125" swimtime="00:01:02.30" />
                    <SPLIT distance="150" swimtime="00:01:16.82" />
                    <SPLIT distance="175" swimtime="00:01:31.95" />
                    <SPLIT distance="200" swimtime="00:01:47.39" />
                    <SPLIT distance="225" swimtime="00:01:57.65" />
                    <SPLIT distance="250" swimtime="00:02:10.42" />
                    <SPLIT distance="275" swimtime="00:02:23.30" />
                    <SPLIT distance="300" swimtime="00:02:36.51" />
                    <SPLIT distance="325" swimtime="00:02:46.97" />
                    <SPLIT distance="350" swimtime="00:02:58.91" />
                    <SPLIT distance="375" swimtime="00:03:11.34" />
                    <SPLIT distance="400" swimtime="00:03:23.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183481" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="105614" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="197514" reactiontime="+22" />
                    <RELAYPOSITION number="4" athleteid="150412" reactiontime="+22" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="United States of America">
              <RESULTS>
                <RESULT eventid="132" place="1" lane="4" heat="1" swimtime="00:06:44.12" reactiontime="+68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.92" />
                    <SPLIT distance="50" swimtime="00:00:23.22" />
                    <SPLIT distance="75" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:00:48.48" />
                    <SPLIT distance="125" swimtime="00:01:01.42" />
                    <SPLIT distance="150" swimtime="00:01:14.47" />
                    <SPLIT distance="175" swimtime="00:01:27.94" />
                    <SPLIT distance="200" swimtime="00:01:41.04" />
                    <SPLIT distance="225" swimtime="00:01:51.94" />
                    <SPLIT distance="250" swimtime="00:02:04.23" />
                    <SPLIT distance="275" swimtime="00:02:16.87" />
                    <SPLIT distance="300" swimtime="00:02:29.59" />
                    <SPLIT distance="325" swimtime="00:02:42.35" />
                    <SPLIT distance="350" swimtime="00:02:55.36" />
                    <SPLIT distance="375" swimtime="00:03:08.51" />
                    <SPLIT distance="400" swimtime="00:03:21.52" />
                    <SPLIT distance="425" swimtime="00:03:32.05" />
                    <SPLIT distance="450" swimtime="00:03:44.49" />
                    <SPLIT distance="475" swimtime="00:03:57.24" />
                    <SPLIT distance="500" swimtime="00:04:10.05" />
                    <SPLIT distance="525" swimtime="00:04:23.13" />
                    <SPLIT distance="550" swimtime="00:04:36.28" />
                    <SPLIT distance="575" swimtime="00:04:49.76" />
                    <SPLIT distance="600" swimtime="00:05:02.96" />
                    <SPLIT distance="625" swimtime="00:05:13.65" />
                    <SPLIT distance="650" swimtime="00:05:25.97" />
                    <SPLIT distance="675" swimtime="00:05:38.48" />
                    <SPLIT distance="700" swimtime="00:05:51.42" />
                    <SPLIT distance="725" swimtime="00:06:04.42" />
                    <SPLIT distance="750" swimtime="00:06:17.69" />
                    <SPLIT distance="775" swimtime="00:06:30.93" />
                    <SPLIT distance="800" swimtime="00:06:44.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150418" reactiontime="+68" />
                    <RELAYPOSITION number="2" athleteid="150412" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="197514" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="145806" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="32" place="1" lane="4" heat="2" swimtime="00:06:53.63" reactiontime="+64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.43" />
                    <SPLIT distance="50" swimtime="00:00:24.28" />
                    <SPLIT distance="75" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:00:50.01" />
                    <SPLIT distance="125" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:16.29" />
                    <SPLIT distance="175" swimtime="00:01:29.78" />
                    <SPLIT distance="200" swimtime="00:01:43.13" />
                    <SPLIT distance="225" swimtime="00:01:53.96" />
                    <SPLIT distance="250" swimtime="00:02:06.81" />
                    <SPLIT distance="275" swimtime="00:02:20.06" />
                    <SPLIT distance="300" swimtime="00:02:33.26" />
                    <SPLIT distance="325" swimtime="00:02:46.48" />
                    <SPLIT distance="350" swimtime="00:02:59.77" />
                    <SPLIT distance="375" swimtime="00:03:13.24" />
                    <SPLIT distance="400" swimtime="00:03:26.37" />
                    <SPLIT distance="425" swimtime="00:03:37.40" />
                    <SPLIT distance="450" swimtime="00:03:50.08" />
                    <SPLIT distance="475" swimtime="00:04:03.25" />
                    <SPLIT distance="500" swimtime="00:04:16.71" />
                    <SPLIT distance="525" swimtime="00:04:30.21" />
                    <SPLIT distance="550" swimtime="00:04:44.01" />
                    <SPLIT distance="575" swimtime="00:04:57.87" />
                    <SPLIT distance="600" swimtime="00:05:11.66" />
                    <SPLIT distance="625" swimtime="00:05:22.53" />
                    <SPLIT distance="650" swimtime="00:05:35.19" />
                    <SPLIT distance="675" swimtime="00:05:48.06" />
                    <SPLIT distance="700" swimtime="00:06:01.01" />
                    <SPLIT distance="725" swimtime="00:06:13.96" />
                    <SPLIT distance="750" swimtime="00:06:27.15" />
                    <SPLIT distance="775" swimtime="00:06:40.45" />
                    <SPLIT distance="800" swimtime="00:06:53.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197514" reactiontime="+64" />
                    <RELAYPOSITION number="2" athleteid="183501" reactiontime="+11" />
                    <RELAYPOSITION number="3" athleteid="214519" reactiontime="+37" />
                    <RELAYPOSITION number="4" athleteid="145806" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="United States of America">
              <RESULTS>
                <RESULT eventid="126" place="5" lane="5" heat="1" swimtime="00:01:24.03" reactiontime="+59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.16" />
                    <SPLIT distance="50" swimtime="00:00:21.16" />
                    <SPLIT distance="75" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:00:41.99" />
                    <SPLIT distance="125" swimtime="00:00:51.93" />
                    <SPLIT distance="150" swimtime="00:01:02.93" />
                    <SPLIT distance="175" swimtime="00:01:12.80" />
                    <SPLIT distance="200" swimtime="00:01:24.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183484" reactiontime="+59" />
                    <RELAYPOSITION number="2" athleteid="197510" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="183481" reactiontime="+26" />
                    <RELAYPOSITION number="4" athleteid="145806" reactiontime="+21" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="26" place="2" lane="5" heat="2" swimtime="00:01:24.07" reactiontime="+62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.22" />
                    <SPLIT distance="50" swimtime="00:00:21.34" />
                    <SPLIT distance="75" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:00:42.29" />
                    <SPLIT distance="125" swimtime="00:00:52.25" />
                    <SPLIT distance="150" swimtime="00:01:03.23" />
                    <SPLIT distance="175" swimtime="00:01:13.13" />
                    <SPLIT distance="200" swimtime="00:01:24.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183484" reactiontime="+62" />
                    <RELAYPOSITION number="2" athleteid="145806" reactiontime="+22" />
                    <RELAYPOSITION number="3" athleteid="183481" reactiontime="+22" />
                    <RELAYPOSITION number="4" athleteid="197510" reactiontime="+40" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="United States of America">
              <RESULTS>
                <RESULT eventid="127" place="4" lane="6" heat="1" swimtime="00:01:29.18" reactiontime="+67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:09.94" />
                    <SPLIT distance="50" swimtime="00:00:20.81" />
                    <SPLIT distance="75" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:00:41.70" />
                    <SPLIT distance="125" swimtime="00:00:52.88" />
                    <SPLIT distance="150" swimtime="00:01:05.23" />
                    <SPLIT distance="175" swimtime="00:01:16.66" />
                    <SPLIT distance="200" swimtime="00:01:29.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124916" reactiontime="+67" />
                    <RELAYPOSITION number="2" athleteid="183484" reactiontime="+33" />
                    <RELAYPOSITION number="3" athleteid="124845" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="150328" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="27" place="4" lane="4" heat="2" swimtime="00:01:29.97" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.29" />
                    <SPLIT distance="50" swimtime="00:00:21.37" />
                    <SPLIT distance="75" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:00:42.18" />
                    <SPLIT distance="125" swimtime="00:00:53.49" />
                    <SPLIT distance="150" swimtime="00:01:06.24" />
                    <SPLIT distance="175" swimtime="00:01:17.48" />
                    <SPLIT distance="200" swimtime="00:01:29.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197510" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="183481" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="202573" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="150328" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="United States of America">
              <RESULTS>
                <RESULT eventid="108" place="2" lane="6" heat="1" swimtime="00:03:26.29" reactiontime="+61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.44" />
                    <SPLIT distance="50" swimtime="00:00:24.38" />
                    <SPLIT distance="75" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:00:51.73" />
                    <SPLIT distance="125" swimtime="00:01:03.15" />
                    <SPLIT distance="150" swimtime="00:01:16.28" />
                    <SPLIT distance="175" swimtime="00:01:29.63" />
                    <SPLIT distance="200" swimtime="00:01:42.90" />
                    <SPLIT distance="225" swimtime="00:01:54.31" />
                    <SPLIT distance="250" swimtime="00:02:07.32" />
                    <SPLIT distance="275" swimtime="00:02:20.76" />
                    <SPLIT distance="300" swimtime="00:02:34.49" />
                    <SPLIT distance="325" swimtime="00:02:45.92" />
                    <SPLIT distance="350" swimtime="00:02:58.97" />
                    <SPLIT distance="375" swimtime="00:03:12.61" />
                    <SPLIT distance="400" swimtime="00:03:26.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183578" reactiontime="+61" />
                    <RELAYPOSITION number="2" athleteid="150313" reactiontime="+34" />
                    <RELAYPOSITION number="3" athleteid="183566" reactiontime="+23" />
                    <RELAYPOSITION number="4" athleteid="124845" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="8" place="4" lane="4" heat="1" swimtime="00:03:31.11" reactiontime="+65">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.15" />
                    <SPLIT distance="50" swimtime="00:00:25.34" />
                    <SPLIT distance="75" swimtime="00:00:39.24" />
                    <SPLIT distance="100" swimtime="00:00:52.83" />
                    <SPLIT distance="125" swimtime="00:01:04.39" />
                    <SPLIT distance="150" swimtime="00:01:17.79" />
                    <SPLIT distance="175" swimtime="00:01:31.85" />
                    <SPLIT distance="200" swimtime="00:01:45.67" />
                    <SPLIT distance="225" swimtime="00:01:57.35" />
                    <SPLIT distance="250" swimtime="00:02:10.63" />
                    <SPLIT distance="275" swimtime="00:02:24.41" />
                    <SPLIT distance="300" swimtime="00:02:38.37" />
                    <SPLIT distance="325" swimtime="00:02:49.77" />
                    <SPLIT distance="350" swimtime="00:03:03.05" />
                    <SPLIT distance="375" swimtime="00:03:17.00" />
                    <SPLIT distance="400" swimtime="00:03:31.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124845" reactiontime="+65" />
                    <RELAYPOSITION number="2" athleteid="183572" reactiontime="+20" />
                    <RELAYPOSITION number="3" athleteid="202573" reactiontime="+38" />
                    <RELAYPOSITION number="4" athleteid="183578" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="United States of America">
              <RESULTS>
                <RESULT eventid="147" place="1" lane="4" heat="1" swimtime="00:03:44.35" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.10" />
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="75" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:00:56.47" />
                    <SPLIT distance="125" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:25.51" />
                    <SPLIT distance="175" swimtime="00:01:42.38" />
                    <SPLIT distance="200" swimtime="00:01:59.35" />
                    <SPLIT distance="225" swimtime="00:02:10.48" />
                    <SPLIT distance="250" swimtime="00:02:24.27" />
                    <SPLIT distance="275" swimtime="00:02:38.82" />
                    <SPLIT distance="300" swimtime="00:02:53.88" />
                    <SPLIT distance="325" swimtime="00:03:04.94" />
                    <SPLIT distance="350" swimtime="00:03:17.85" />
                    <SPLIT distance="375" swimtime="00:03:31.16" />
                    <SPLIT distance="400" swimtime="00:03:44.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183566" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="130153" reactiontime="+38" />
                    <RELAYPOSITION number="3" athleteid="183578" reactiontime="+27" />
                    <RELAYPOSITION number="4" athleteid="150313" reactiontime="+31" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="47" place="1" lane="5" heat="1" swimtime="00:03:47.67" reactiontime="+70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                    <SPLIT distance="75" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:00:56.60" />
                    <SPLIT distance="125" swimtime="00:01:10.02" />
                    <SPLIT distance="150" swimtime="00:01:26.30" />
                    <SPLIT distance="175" swimtime="00:01:43.31" />
                    <SPLIT distance="200" swimtime="00:02:00.63" />
                    <SPLIT distance="225" swimtime="00:02:11.85" />
                    <SPLIT distance="250" swimtime="00:02:25.83" />
                    <SPLIT distance="275" swimtime="00:02:40.33" />
                    <SPLIT distance="300" swimtime="00:02:55.09" />
                    <SPLIT distance="325" swimtime="00:03:06.88" />
                    <SPLIT distance="350" swimtime="00:03:20.18" />
                    <SPLIT distance="375" swimtime="00:03:34.05" />
                    <SPLIT distance="400" swimtime="00:03:47.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150328" reactiontime="+70" />
                    <RELAYPOSITION number="2" athleteid="130153" reactiontime="+29" />
                    <RELAYPOSITION number="3" athleteid="150313" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="124845" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="United States of America">
              <RESULTS>
                <RESULT eventid="117" place="3" lane="4" heat="1" swimtime="00:07:34.70" reactiontime="+74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="75" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:00:55.39" />
                    <SPLIT distance="125" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:24.64" />
                    <SPLIT distance="175" swimtime="00:01:39.51" />
                    <SPLIT distance="200" swimtime="00:01:53.90" />
                    <SPLIT distance="225" swimtime="00:02:06.24" />
                    <SPLIT distance="250" swimtime="00:02:20.45" />
                    <SPLIT distance="275" swimtime="00:02:34.80" />
                    <SPLIT distance="300" swimtime="00:02:49.24" />
                    <SPLIT distance="325" swimtime="00:03:03.80" />
                    <SPLIT distance="350" swimtime="00:03:18.33" />
                    <SPLIT distance="375" swimtime="00:03:33.12" />
                    <SPLIT distance="400" swimtime="00:03:47.38" />
                    <SPLIT distance="425" swimtime="00:03:59.17" />
                    <SPLIT distance="450" swimtime="00:04:12.70" />
                    <SPLIT distance="475" swimtime="00:04:26.86" />
                    <SPLIT distance="500" swimtime="00:04:41.15" />
                    <SPLIT distance="525" swimtime="00:04:55.53" />
                    <SPLIT distance="550" swimtime="00:05:10.26" />
                    <SPLIT distance="575" swimtime="00:05:25.20" />
                    <SPLIT distance="600" swimtime="00:05:39.61" />
                    <SPLIT distance="625" swimtime="00:05:51.98" />
                    <SPLIT distance="650" swimtime="00:06:06.05" />
                    <SPLIT distance="675" swimtime="00:06:20.57" />
                    <SPLIT distance="700" swimtime="00:06:35.39" />
                    <SPLIT distance="725" swimtime="00:06:50.18" />
                    <SPLIT distance="750" swimtime="00:07:05.14" />
                    <SPLIT distance="775" swimtime="00:07:20.21" />
                    <SPLIT distance="800" swimtime="00:07:34.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150328" reactiontime="+74" />
                    <RELAYPOSITION number="2" athleteid="143364" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="183572" reactiontime="+18" />
                    <RELAYPOSITION number="4" athleteid="105648" reactiontime="+24" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="17" place="1" lane="4" heat="1" swimtime="00:07:42.91" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.91" />
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="75" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:00:56.86" />
                    <SPLIT distance="125" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:26.97" />
                    <SPLIT distance="175" swimtime="00:01:41.99" />
                    <SPLIT distance="200" swimtime="00:01:56.61" />
                    <SPLIT distance="225" swimtime="00:02:09.09" />
                    <SPLIT distance="250" swimtime="00:02:23.33" />
                    <SPLIT distance="275" swimtime="00:02:37.68" />
                    <SPLIT distance="300" swimtime="00:02:52.18" />
                    <SPLIT distance="325" swimtime="00:03:06.88" />
                    <SPLIT distance="350" swimtime="00:03:21.65" />
                    <SPLIT distance="375" swimtime="00:03:36.49" />
                    <SPLIT distance="400" swimtime="00:03:51.00" />
                    <SPLIT distance="425" swimtime="00:04:03.47" />
                    <SPLIT distance="450" swimtime="00:04:17.61" />
                    <SPLIT distance="475" swimtime="00:04:32.07" />
                    <SPLIT distance="500" swimtime="00:04:46.99" />
                    <SPLIT distance="525" swimtime="00:05:01.90" />
                    <SPLIT distance="550" swimtime="00:05:17.05" />
                    <SPLIT distance="575" swimtime="00:05:32.23" />
                    <SPLIT distance="600" swimtime="00:05:47.03" />
                    <SPLIT distance="625" swimtime="00:05:59.67" />
                    <SPLIT distance="650" swimtime="00:06:14.07" />
                    <SPLIT distance="675" swimtime="00:06:28.64" />
                    <SPLIT distance="700" swimtime="00:06:43.50" />
                    <SPLIT distance="725" swimtime="00:06:58.41" />
                    <SPLIT distance="750" swimtime="00:07:13.45" />
                    <SPLIT distance="775" swimtime="00:07:28.36" />
                    <SPLIT distance="800" swimtime="00:07:42.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124845" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="143364" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="213247" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="105648" reactiontime="+30" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="United States of America">
              <RESULTS>
                <RESULT eventid="125" place="1" lane="3" heat="1" swimtime="00:01:33.89" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.42" />
                    <SPLIT distance="50" swimtime="00:00:24.08" />
                    <SPLIT distance="75" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:00:47.38" />
                    <SPLIT distance="125" swimtime="00:00:58.82" />
                    <SPLIT distance="150" swimtime="00:01:11.12" />
                    <SPLIT distance="175" swimtime="00:01:21.94" />
                    <SPLIT distance="200" swimtime="00:01:33.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183578" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="183566" reactiontime="+4" />
                    <RELAYPOSITION number="3" athleteid="124845" reactiontime="+36" />
                    <RELAYPOSITION number="4" athleteid="150313" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="25" place="3" lane="4" heat="2" swimtime="00:01:36.17" reactiontime="+63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.82" />
                    <SPLIT distance="50" swimtime="00:00:24.16" />
                    <SPLIT distance="75" swimtime="00:00:35.77" />
                    <SPLIT distance="100" swimtime="00:00:48.50" />
                    <SPLIT distance="125" swimtime="00:00:59.69" />
                    <SPLIT distance="150" swimtime="00:01:12.42" />
                    <SPLIT distance="175" swimtime="00:01:23.69" />
                    <SPLIT distance="200" swimtime="00:01:36.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="124845" reactiontime="+63" />
                    <RELAYPOSITION number="2" athleteid="183572" reactiontime="+13" />
                    <RELAYPOSITION number="3" athleteid="202573" reactiontime="+29" />
                    <RELAYPOSITION number="4" athleteid="150328" reactiontime="+23" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="United States of America">
              <RESULTS>
                <RESULT eventid="134" place="2" lane="1" heat="1" swimtime="00:01:42.41" reactiontime="+58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.64" />
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                    <SPLIT distance="75" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:00:54.75" />
                    <SPLIT distance="125" swimtime="00:01:06.00" />
                    <SPLIT distance="150" swimtime="00:01:19.69" />
                    <SPLIT distance="175" swimtime="00:01:30.38" />
                    <SPLIT distance="200" swimtime="00:01:42.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183566" reactiontime="+58" />
                    <RELAYPOSITION number="2" athleteid="130153" reactiontime="+24" />
                    <RELAYPOSITION number="3" athleteid="183578" reactiontime="+38" />
                    <RELAYPOSITION number="4" athleteid="150313" reactiontime="+25" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="34" place="7" lane="4" heat="1" swimtime="00:01:46.58" reactiontime="+73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.70" />
                    <SPLIT distance="50" swimtime="00:00:27.18" />
                    <SPLIT distance="75" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:00:57.32" />
                    <SPLIT distance="125" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:22.49" />
                    <SPLIT distance="175" swimtime="00:01:33.94" />
                    <SPLIT distance="200" swimtime="00:01:46.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="150328" reactiontime="+73" />
                    <RELAYPOSITION number="2" athleteid="156655" reactiontime="+16" />
                    <RELAYPOSITION number="3" athleteid="124845" reactiontime="+34" />
                    <RELAYPOSITION number="4" athleteid="202573" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="United States of America">
              <RESULTS>
                <RESULT eventid="111" place="1" lane="4" heat="1" swimtime="00:01:35.15" reactiontime="+51">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.95" />
                    <SPLIT distance="50" swimtime="00:00:22.37" />
                    <SPLIT distance="75" swimtime="00:00:33.53" />
                    <SPLIT distance="100" swimtime="00:00:47.33" />
                    <SPLIT distance="125" swimtime="00:00:58.10" />
                    <SPLIT distance="150" swimtime="00:01:11.42" />
                    <SPLIT distance="175" swimtime="00:01:22.55" />
                    <SPLIT distance="200" swimtime="00:01:35.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="105644" reactiontime="+51" />
                    <RELAYPOSITION number="2" athleteid="105614" reactiontime="+19" />
                    <RELAYPOSITION number="3" athleteid="150313" reactiontime="+28" />
                    <RELAYPOSITION number="4" athleteid="183578" reactiontime="+35" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="11" place="1" lane="4" heat="2" swimtime="00:01:36.83" reactiontime="+52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.25" />
                    <SPLIT distance="50" swimtime="00:00:22.98" />
                    <SPLIT distance="75" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:00:48.54" />
                    <SPLIT distance="125" swimtime="00:00:59.56" />
                    <SPLIT distance="150" swimtime="00:01:12.91" />
                    <SPLIT distance="175" swimtime="00:01:24.37" />
                    <SPLIT distance="200" swimtime="00:01:36.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="197510" reactiontime="+52" />
                    <RELAYPOSITION number="2" athleteid="124916" reactiontime="+36" />
                    <RELAYPOSITION number="3" athleteid="150313" reactiontime="+35" />
                    <RELAYPOSITION number="4" athleteid="150328" reactiontime="+38" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY number="1" agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="United States of America">
              <RESULTS>
                <RESULT eventid="135" place="2" lane="2" heat="1" swimtime="00:01:30.37" reactiontime="+49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.05" />
                    <SPLIT distance="50" swimtime="00:00:22.61" />
                    <SPLIT distance="75" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:00:47.85" />
                    <SPLIT distance="125" swimtime="00:00:57.71" />
                    <SPLIT distance="150" swimtime="00:01:09.98" />
                    <SPLIT distance="175" swimtime="00:01:19.56" />
                    <SPLIT distance="200" swimtime="00:01:30.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="105644" reactiontime="+49" />
                    <RELAYPOSITION number="2" athleteid="105614" reactiontime="+25" />
                    <RELAYPOSITION number="3" athleteid="197510" reactiontime="+24" />
                    <RELAYPOSITION number="4" athleteid="124916" reactiontime="+37" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="35" place="5" lane="4" heat="2" swimtime="00:01:32.67" reactiontime="+60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.46" />
                    <SPLIT distance="50" swimtime="00:00:23.34" />
                    <SPLIT distance="75" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:00:48.94" />
                    <SPLIT distance="125" swimtime="00:00:59.04" />
                    <SPLIT distance="150" swimtime="00:01:11.33" />
                    <SPLIT distance="175" swimtime="00:01:21.54" />
                    <SPLIT distance="200" swimtime="00:01:32.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="1" athleteid="183481" reactiontime="+60" />
                    <RELAYPOSITION number="2" athleteid="105614" reactiontime="+30" />
                    <RELAYPOSITION number="3" athleteid="197514" reactiontime="+25" />
                    <RELAYPOSITION number="4" athleteid="150418" reactiontime="+32" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB name="Uzbekistan" shortname="UZB" code="UZB" nation="UZB" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="195293" lastname="USMONOV" firstname="Eldor" gender="M" birthdate="2004-01-31">
              <ENTRIES>
                <ENTRY entrytime="00:00:53.54" eventid="39" heat="4" lane="1">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
                <ENTRY entrytime="00:00:24.07" eventid="5" heat="5" lane="8">
                  <MEETINFO date="2022-08-17" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="39" place="32" lane="1" heat="4" heatid="40039" swimtime="00:00:52.19" reactiontime="+66" points="767">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.61" />
                    <SPLIT distance="50" swimtime="00:00:23.82" />
                    <SPLIT distance="75" swimtime="00:00:37.56" />
                    <SPLIT distance="100" swimtime="00:00:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="5" place="45" lane="8" heat="5" heatid="50005" swimtime="00:00:23.50" reactiontime="+75" points="792">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.63" />
                    <SPLIT distance="50" swimtime="00:00:23.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106908" lastname="TARASENKO" firstname="Aleksey" gender="M" birthdate="1999-05-13">
              <ENTRIES>
                <ENTRY entrytime="00:00:48.45" eventid="14" heat="7" lane="8">
                  <MEETINFO date="2021-12-20" />
                </ENTRY>
                <ENTRY entrytime="00:00:21.91" eventid="31" heat="7" lane="3">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="14" place="38" lane="8" heat="7" heatid="70014" swimtime="00:00:47.82" reactiontime="+65" points="824">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.96" />
                    <SPLIT distance="50" swimtime="00:00:23.18" />
                    <SPLIT distance="75" swimtime="00:00:35.46" />
                    <SPLIT distance="100" swimtime="00:00:47.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="31" place="36" lane="3" heat="7" heatid="70031" swimtime="00:00:21.59" reactiontime="+61" points="814">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:10.40" />
                    <SPLIT distance="50" swimtime="00:00:21.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB name="Zimbabwe" shortname="ZIM" code="ZIM" nation="ZIM" type="NOC">
          <ATHLETES>
            <ATHLETE athleteid="129273" lastname="O'HARA" firstname="Liam" gender="M" birthdate="2001-02-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.01" eventid="16" heat="2" lane="4">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="00:02:07.12" eventid="7" heat="1" lane="5">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="16" place="48" lane="4" heat="2" heatid="20016" swimtime="00:01:01.31" reactiontime="+61" points="733">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.98" />
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="75" swimtime="00:00:44.62" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="7" place="35" lane="5" heat="1" heatid="10007" swimtime="00:02:04.90" reactiontime="+65" points="676">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.07" />
                    <SPLIT distance="50" swimtime="00:00:26.99" />
                    <SPLIT distance="75" swimtime="00:00:43.48" />
                    <SPLIT distance="100" swimtime="00:00:58.98" />
                    <SPLIT distance="125" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:01:33.57" />
                    <SPLIT distance="175" swimtime="00:01:49.80" />
                    <SPLIT distance="200" swimtime="00:02:04.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="106974" lastname="DAVIS" firstname="Liam" gender="M" birthdate="2000-04-04">
              <ENTRIES>
                <ENTRY entrytime="00:02:15.28" eventid="29" heat="1" lane="5">
                  <MEETINFO date="2021-12-18" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="29" place="29" lane="5" heat="1" heatid="10029" swimtime="00:02:13.99" reactiontime="+67" points="721">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.13" />
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="75" swimtime="00:00:47.02" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="125" swimtime="00:01:20.97" />
                    <SPLIT distance="150" swimtime="00:01:38.31" />
                    <SPLIT distance="175" swimtime="00:01:56.02" />
                    <SPLIT distance="200" swimtime="00:02:13.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="168820" lastname="KATAI" firstname="Donata" gender="F" birthdate="2004-05-07">
              <ENTRIES>
                <ENTRY entrytime="00:01:02.73" eventid="2" heat="2" lane="4">
                  <MEETINFO date="2021-07-25" />
                </ENTRY>
                <ENTRY entrytime="00:00:29.81" eventid="18" heat="3" lane="5">
                  <MEETINFO date="2022-06-21" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="2" place="37" lane="4" heat="2" heatid="20002" swimtime="00:01:01.85" reactiontime="+61" points="698">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.54" />
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="75" swimtime="00:00:46.25" />
                    <SPLIT distance="100" swimtime="00:01:01.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="18" place="35" lane="5" heat="3" heatid="30018" swimtime="00:00:28.83" reactiontime="+60" points="673">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.21" />
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE athleteid="201959" lastname="MJIMBA" firstname="Nomvula" gender="F" birthdate="2002-03-17">
              <ENTRIES>
                <ENTRY entrytime="00:01:00.32" eventid="13" heat="4" lane="8">
                  <MEETINFO date="2022-08-11" />
                </ENTRY>
                <ENTRY entrytime="00:00:27.81" eventid="30" heat="4" lane="8">
                  <MEETINFO date="2022-08-13" />
                </ENTRY>
              </ENTRIES>
              <RESULTS>
                <RESULT eventid="13" place="51" lane="8" heat="4" heatid="40013" swimtime="00:00:59.81" reactiontime="+63" points="593">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.55" />
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="75" swimtime="00:00:44.09" />
                    <SPLIT distance="100" swimtime="00:00:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="30" place="39" lane="8" heat="4" heatid="40030" swimtime="00:00:27.15" reactiontime="+60" points="602">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.09" />
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>