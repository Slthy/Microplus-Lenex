<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Schwimmclub Aarefisch" version="11.75236">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Aarau" name="Aargau Open 2022" course="SCM" deadline="2022-11-25" entrytype="OPEN" hostclub="Schwimmclub Aarefisch, Aarau" hostclub.url="http://www.aarefisch.ch" organizer="Schwimmclub Aarefisch, Aarau" organizer.url="http://www.aarefisch.ch" reservecount="2" result.url="https://live.swimrankings.net/32190/" startmethod="1" timing="AUTOMATIC" type="SUI.IM" state="AG" nation="SUI">
      <AGEDATE value="2022-12-05" type="YEAR" />
      <POOL name="Hallenbad Telli Aarau" lanemin="1" lanemax="4" />
      <FACILITY city="Aarau" name="Hallenbad Telli Aarau" nation="SUI" state="AG" street="Tellistrasse 80" zip="5000" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <CONTACT city="Aarau" email="wettkaempfe@aarefisch.ch" name="Schwimmclub Aarefisch, Aarau" street="Geschäftsstelle " street2="Weihermattstrasse 74/76" zip="5000" />
      <SESSIONS>
        <SESSION date="2022-12-03" daytime="08:30" name="De / Rü Vormittag" number="1" officialmeeting="08:00" teamleadermeeting="07:30" warmupfrom="07:15" warmupuntil="08:20">
          <EVENTS>
            <EVENT eventid="1064" daytime="08:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1065" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13079" />
                    <RANKING order="2" place="2" resultid="13017" />
                    <RANKING order="3" place="3" resultid="12957" />
                    <RANKING order="4" place="4" resultid="14121" />
                    <RANKING order="5" place="5" resultid="12721" />
                    <RANKING order="6" place="6" resultid="14235" />
                    <RANKING order="7" place="7" resultid="13900" />
                    <RANKING order="8" place="8" resultid="13999" />
                    <RANKING order="9" place="9" resultid="14441" />
                    <RANKING order="10" place="10" resultid="14424" />
                    <RANKING order="11" place="-1" resultid="14384" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14513" daytime="08:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14514" daytime="08:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14515" daytime="08:33" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="08:35" gender="M" number="2" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1137" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13030" />
                    <RANKING order="2" place="2" resultid="14028" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14516" daytime="08:35" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="08:37" gender="F" number="3" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12781" />
                    <RANKING order="2" place="2" resultid="12134" />
                    <RANKING order="3" place="3" resultid="12709" />
                    <RANKING order="4" place="4" resultid="12883" />
                    <RANKING order="5" place="5" resultid="12786" />
                    <RANKING order="6" place="6" resultid="14023" />
                    <RANKING order="7" place="7" resultid="12500" />
                    <RANKING order="8" place="8" resultid="14060" />
                    <RANKING order="9" place="9" resultid="14380" />
                    <RANKING order="10" place="10" resultid="14350" />
                    <RANKING order="11" place="11" resultid="14213" />
                    <RANKING order="12" place="-1" resultid="14103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12697" />
                    <RANKING order="2" place="2" resultid="12684" />
                    <RANKING order="3" place="-1" resultid="12146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12702" />
                    <RANKING order="2" place="2" resultid="14240" />
                    <RANKING order="3" place="3" resultid="13198" />
                    <RANKING order="4" place="4" resultid="12743" />
                    <RANKING order="5" place="5" resultid="14033" />
                    <RANKING order="6" place="6" resultid="12813" />
                    <RANKING order="7" place="7" resultid="12545" />
                    <RANKING order="8" place="8" resultid="12573" />
                    <RANKING order="9" place="-1" resultid="13970" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14517" daytime="08:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14518" daytime="08:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14519" daytime="08:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14520" daytime="08:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14521" daytime="08:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14522" daytime="08:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="08:51" gender="M" number="4" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1155" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13074" />
                    <RANKING order="2" place="2" resultid="14051" />
                    <RANKING order="3" place="3" resultid="12791" />
                    <RANKING order="4" place="4" resultid="14098" />
                    <RANKING order="5" place="5" resultid="12535" />
                    <RANKING order="6" place="6" resultid="12568" />
                    <RANKING order="7" place="-1" resultid="13134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="13848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12966" />
                    <RANKING order="2" place="2" resultid="14169" />
                    <RANKING order="3" place="3" resultid="12808" />
                    <RANKING order="4" place="4" resultid="12712" />
                    <RANKING order="5" place="5" resultid="12768" />
                    <RANKING order="6" place="6" resultid="12726" />
                    <RANKING order="7" place="7" resultid="14164" />
                    <RANKING order="8" place="-1" resultid="12558" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14523" daytime="08:51" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14524" daytime="08:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14525" daytime="08:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14526" daytime="08:59" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="09:01" gender="F" number="5" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14820" />
                    <RANKING order="2" place="2" resultid="13870" />
                    <RANKING order="3" place="3" resultid="13852" />
                    <RANKING order="4" place="4" resultid="14226" />
                    <RANKING order="5" place="4" resultid="14396" />
                    <RANKING order="6" place="6" resultid="14015" />
                    <RANKING order="7" place="7" resultid="12607" />
                    <RANKING order="8" place="8" resultid="13912" />
                    <RANKING order="9" place="9" resultid="14149" />
                    <RANKING order="10" place="-1" resultid="12662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13080" />
                    <RANKING order="2" place="2" resultid="14122" />
                    <RANKING order="3" place="3" resultid="13018" />
                    <RANKING order="4" place="4" resultid="12722" />
                    <RANKING order="5" place="5" resultid="12958" />
                    <RANKING order="6" place="6" resultid="14236" />
                    <RANKING order="7" place="7" resultid="14421" />
                    <RANKING order="8" place="8" resultid="13376" />
                    <RANKING order="9" place="9" resultid="14133" />
                    <RANKING order="10" place="10" resultid="14000" />
                    <RANKING order="11" place="11" resultid="14438" />
                    <RANKING order="12" place="12" resultid="13966" />
                    <RANKING order="13" place="13" resultid="14047" />
                    <RANKING order="14" place="14" resultid="14272" />
                    <RANKING order="15" place="-1" resultid="14385" />
                    <RANKING order="16" place="-1" resultid="13901" />
                    <RANKING order="17" place="-1" resultid="14343" />
                    <RANKING order="18" place="-1" resultid="12630" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14527" daytime="09:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14528" daytime="09:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14529" daytime="09:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14530" daytime="09:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14531" daytime="09:07" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14532" daytime="09:09" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14533" daytime="09:10" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:12" gender="M" number="6" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1143" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12773" />
                    <RANKING order="2" place="2" resultid="14082" />
                    <RANKING order="3" place="3" resultid="12778" />
                    <RANKING order="4" place="4" resultid="14157" />
                    <RANKING order="5" place="5" resultid="14126" />
                    <RANKING order="6" place="6" resultid="14258" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14029" />
                    <RANKING order="2" place="2" resultid="13031" />
                    <RANKING order="3" place="3" resultid="14511" />
                    <RANKING order="4" place="4" resultid="14069" />
                    <RANKING order="5" place="5" resultid="14043" />
                    <RANKING order="6" place="6" resultid="14403" />
                    <RANKING order="7" place="7" resultid="14335" />
                    <RANKING order="8" place="-1" resultid="12693" />
                    <RANKING order="9" place="-1" resultid="13856" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14534" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14535" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14536" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14537" daytime="09:17" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1078" daytime="09:19" gender="F" number="7" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1176" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14339" />
                    <RANKING order="2" place="2" resultid="12782" />
                    <RANKING order="3" place="3" resultid="12884" />
                    <RANKING order="4" place="4" resultid="12118" />
                    <RANKING order="5" place="5" resultid="14024" />
                    <RANKING order="6" place="6" resultid="14061" />
                    <RANKING order="7" place="7" resultid="14381" />
                    <RANKING order="8" place="8" resultid="12748" />
                    <RANKING order="9" place="9" resultid="12787" />
                    <RANKING order="10" place="10" resultid="13013" />
                    <RANKING order="11" place="11" resultid="12710" />
                    <RANKING order="12" place="12" resultid="14214" />
                    <RANKING order="13" place="13" resultid="12501" />
                    <RANKING order="14" place="14" resultid="12913" />
                    <RANKING order="15" place="15" resultid="13808" />
                    <RANKING order="16" place="16" resultid="12114" />
                    <RANKING order="17" place="17" resultid="12800" />
                    <RANKING order="18" place="18" resultid="13147" />
                    <RANKING order="19" place="19" resultid="13915" />
                    <RANKING order="20" place="20" resultid="14369" />
                    <RANKING order="21" place="21" resultid="12804" />
                    <RANKING order="22" place="22" resultid="14359" />
                    <RANKING order="23" place="-1" resultid="13310" />
                    <RANKING order="24" place="-1" resultid="14392" />
                    <RANKING order="25" place="-1" resultid="12488" />
                    <RANKING order="26" place="-1" resultid="12756" />
                    <RANKING order="27" place="-1" resultid="12899" />
                    <RANKING order="28" place="-1" resultid="13089" />
                    <RANKING order="29" place="-1" resultid="13874" />
                    <RANKING order="30" place="-1" resultid="13888" />
                    <RANKING order="31" place="-1" resultid="13919" />
                    <RANKING order="32" place="-1" resultid="14104" />
                    <RANKING order="33" place="-1" resultid="14372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12685" />
                    <RANKING order="2" place="2" resultid="13839" />
                    <RANKING order="3" place="3" resultid="13928" />
                    <RANKING order="4" place="4" resultid="13896" />
                    <RANKING order="5" place="5" resultid="12698" />
                    <RANKING order="6" place="6" resultid="14376" />
                    <RANKING order="7" place="7" resultid="13308" />
                    <RANKING order="8" place="8" resultid="12975" />
                    <RANKING order="9" place="9" resultid="12531" />
                    <RANKING order="10" place="10" resultid="14245" />
                    <RANKING order="11" place="11" resultid="14019" />
                    <RANKING order="12" place="12" resultid="12669" />
                    <RANKING order="13" place="13" resultid="13105" />
                    <RANKING order="14" place="14" resultid="12505" />
                    <RANKING order="15" place="-1" resultid="12689" />
                    <RANKING order="16" place="-1" resultid="13005" />
                    <RANKING order="17" place="-1" resultid="13043" />
                    <RANKING order="18" place="-1" resultid="13155" />
                    <RANKING order="19" place="-1" resultid="13293" />
                    <RANKING order="20" place="-1" resultid="12509" />
                    <RANKING order="21" place="-1" resultid="13026" />
                    <RANKING order="22" place="-1" resultid="12147" />
                    <RANKING order="23" place="-1" resultid="12619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12703" />
                    <RANKING order="2" place="2" resultid="14241" />
                    <RANKING order="3" place="3" resultid="12744" />
                    <RANKING order="4" place="4" resultid="14034" />
                    <RANKING order="5" place="5" resultid="12920" />
                    <RANKING order="6" place="6" resultid="12814" />
                    <RANKING order="7" place="7" resultid="12574" />
                    <RANKING order="8" place="8" resultid="12932" />
                    <RANKING order="9" place="9" resultid="12546" />
                    <RANKING order="10" place="10" resultid="14361" />
                    <RANKING order="11" place="11" resultid="13819" />
                    <RANKING order="12" place="12" resultid="13971" />
                    <RANKING order="13" place="13" resultid="13245" />
                    <RANKING order="14" place="14" resultid="12962" />
                    <RANKING order="15" place="15" resultid="14430" />
                    <RANKING order="16" place="16" resultid="14056" />
                    <RANKING order="17" place="17" resultid="13832" />
                    <RANKING order="18" place="18" resultid="13055" />
                    <RANKING order="19" place="19" resultid="13314" />
                    <RANKING order="20" place="20" resultid="13302" />
                    <RANKING order="21" place="21" resultid="12177" />
                    <RANKING order="22" place="-1" resultid="12891" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14538" daytime="09:19" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14539" daytime="09:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14540" daytime="09:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14541" daytime="09:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14542" daytime="09:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14543" daytime="09:32" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14544" daytime="09:35" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14545" daytime="09:37" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14546" daytime="09:39" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14547" daytime="09:41" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14548" daytime="09:43" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14549" daytime="09:46" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14550" daytime="09:48" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14551" daytime="09:50" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14552" daytime="09:52" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14553" daytime="09:54" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="14554" daytime="09:56" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1081" daytime="10:00" gender="M" number="8" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1162" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12928" />
                    <RANKING order="2" place="2" resultid="12796" />
                    <RANKING order="3" place="3" resultid="14448" />
                    <RANKING order="4" place="4" resultid="14365" />
                    <RANKING order="5" place="5" resultid="12731" />
                    <RANKING order="6" place="6" resultid="13009" />
                    <RANKING order="7" place="7" resultid="14117" />
                    <RANKING order="8" place="8" resultid="14094" />
                    <RANKING order="9" place="9" resultid="13159" />
                    <RANKING order="10" place="10" resultid="14434" />
                    <RANKING order="11" place="11" resultid="12554" />
                    <RANKING order="12" place="12" resultid="12739" />
                    <RANKING order="13" place="13" resultid="13957" />
                    <RANKING order="14" place="14" resultid="13909" />
                    <RANKING order="15" place="15" resultid="14222" />
                    <RANKING order="16" place="16" resultid="14426" />
                    <RANKING order="17" place="17" resultid="12138" />
                    <RANKING order="18" place="18" resultid="13039" />
                    <RANKING order="19" place="19" resultid="13132" />
                    <RANKING order="20" place="20" resultid="13112" />
                    <RANKING order="21" place="21" resultid="12550" />
                    <RANKING order="22" place="-1" resultid="12611" />
                    <RANKING order="23" place="-1" resultid="12603" />
                    <RANKING order="24" place="-1" resultid="13035" />
                    <RANKING order="25" place="-1" resultid="13284" />
                    <RANKING order="26" place="-1" resultid="13849" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14099" />
                    <RANKING order="2" place="2" resultid="12792" />
                    <RANKING order="3" place="3" resultid="14052" />
                    <RANKING order="4" place="4" resultid="13804" />
                    <RANKING order="5" place="5" resultid="12536" />
                    <RANKING order="6" place="6" resultid="12760" />
                    <RANKING order="7" place="7" resultid="13075" />
                    <RANKING order="8" place="8" resultid="12735" />
                    <RANKING order="9" place="9" resultid="12752" />
                    <RANKING order="10" place="10" resultid="12910" />
                    <RANKING order="11" place="11" resultid="14113" />
                    <RANKING order="12" place="12" resultid="13047" />
                    <RANKING order="13" place="13" resultid="13945" />
                    <RANKING order="14" place="14" resultid="14249" />
                    <RANKING order="15" place="-1" resultid="12717" />
                    <RANKING order="16" place="-1" resultid="12569" />
                    <RANKING order="17" place="-1" resultid="14179" />
                    <RANKING order="18" place="-1" resultid="13135" />
                    <RANKING order="19" place="-1" resultid="14400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12967" />
                    <RANKING order="2" place="2" resultid="12809" />
                    <RANKING order="3" place="3" resultid="14170" />
                    <RANKING order="4" place="4" resultid="12713" />
                    <RANKING order="5" place="5" resultid="12903" />
                    <RANKING order="6" place="6" resultid="12863" />
                    <RANKING order="7" place="7" resultid="14165" />
                    <RANKING order="8" place="8" resultid="12727" />
                    <RANKING order="9" place="9" resultid="13260" />
                    <RANKING order="10" place="10" resultid="12895" />
                    <RANKING order="11" place="11" resultid="12769" />
                    <RANKING order="12" place="12" resultid="14065" />
                    <RANKING order="13" place="13" resultid="12169" />
                    <RANKING order="14" place="14" resultid="13369" />
                    <RANKING order="15" place="15" resultid="12559" />
                    <RANKING order="16" place="16" resultid="12764" />
                    <RANKING order="17" place="17" resultid="13815" />
                    <RANKING order="18" place="18" resultid="12638" />
                    <RANKING order="19" place="19" resultid="13953" />
                    <RANKING order="20" place="20" resultid="14153" />
                    <RANKING order="21" place="21" resultid="13942" />
                    <RANKING order="22" place="-1" resultid="13051" />
                    <RANKING order="23" place="-1" resultid="13063" />
                    <RANKING order="24" place="-1" resultid="13365" />
                    <RANKING order="25" place="-1" resultid="13387" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14558" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14559" daytime="10:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14560" daytime="10:07" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14561" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14562" daytime="10:12" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14563" daytime="10:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14564" daytime="10:17" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14565" daytime="10:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14566" daytime="10:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14567" daytime="10:24" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14568" daytime="10:27" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14569" daytime="10:29" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14570" daytime="10:31" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14571" daytime="10:33" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14572" daytime="10:35" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14573" daytime="10:37" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2022-12-03" daytime="10:45" name="Staffeln Freistil Vormittag" number="2">
          <EVENTS>
            <EVENT eventid="1084" daytime="10:45" gender="F" number="9" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="CHF" value="1800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1085" agemax="12" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12821" />
                    <RANKING order="2" place="2" resultid="14809" />
                    <RANKING order="3" place="3" resultid="12937" />
                    <RANKING order="4" place="4" resultid="14457" />
                    <RANKING order="5" place="5" resultid="13171" />
                    <RANKING order="6" place="6" resultid="13335" />
                    <RANKING order="7" place="7" resultid="12822" />
                    <RANKING order="8" place="8" resultid="12578" />
                    <RANKING order="9" place="9" resultid="13842" />
                    <RANKING order="10" place="10" resultid="13977" />
                    <RANKING order="11" place="11" resultid="14810" />
                    <RANKING order="12" place="12" resultid="14459" />
                    <RANKING order="13" place="13" resultid="12823" />
                    <RANKING order="14" place="14" resultid="13337" />
                    <RANKING order="15" place="15" resultid="13175" />
                    <RANKING order="16" place="16" resultid="14811" />
                    <RANKING order="17" place="17" resultid="13978" />
                    <RANKING order="18" place="18" resultid="12580" />
                    <RANKING order="19" place="19" resultid="14812" />
                    <RANKING order="20" place="-1" resultid="12190" />
                    <RANKING order="21" place="-1" resultid="13173" />
                    <RANKING order="22" place="-1" resultid="14460" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14576" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14577" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14578" daytime="10:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14579" daytime="10:57" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14580" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14817" daytime="11:03" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="11:06" gender="M" number="10" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="CHF" value="1800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="12" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12817" />
                    <RANKING order="2" place="2" resultid="14813" />
                    <RANKING order="3" place="3" resultid="12935" />
                    <RANKING order="4" place="4" resultid="14814" />
                    <RANKING order="5" place="5" resultid="13333" />
                    <RANKING order="6" place="6" resultid="12819" />
                    <RANKING order="7" place="7" resultid="12577" />
                    <RANKING order="8" place="8" resultid="14815" />
                    <RANKING order="9" place="9" resultid="13169" />
                    <RANKING order="10" place="10" resultid="13974" />
                    <RANKING order="11" place="11" resultid="14816" />
                    <RANKING order="12" place="-1" resultid="13167" />
                    <RANKING order="13" place="-1" resultid="12818" />
                    <RANKING order="14" place="-1" resultid="14456" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14581" daytime="11:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14582" daytime="11:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14583" daytime="11:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14818" daytime="11:17" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2022-12-03" daytime="11:24" endtime="14:56" name="Br / Cr Vormittag" number="3">
          <EVENTS>
            <EVENT eventid="1088" daytime="11:24" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1145" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14821" />
                    <RANKING order="2" place="2" resultid="14016" />
                    <RANKING order="3" place="3" resultid="13871" />
                    <RANKING order="4" place="4" resultid="14227" />
                    <RANKING order="5" place="5" resultid="12608" />
                    <RANKING order="6" place="6" resultid="13853" />
                    <RANKING order="7" place="7" resultid="14150" />
                    <RANKING order="8" place="-1" resultid="14398" />
                    <RANKING order="9" place="-1" resultid="12663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13081" />
                    <RANKING order="2" place="2" resultid="13019" />
                    <RANKING order="3" place="3" resultid="12723" />
                    <RANKING order="4" place="4" resultid="12959" />
                    <RANKING order="5" place="5" resultid="14123" />
                    <RANKING order="6" place="6" resultid="14387" />
                    <RANKING order="7" place="7" resultid="14001" />
                    <RANKING order="8" place="8" resultid="14237" />
                    <RANKING order="9" place="9" resultid="14048" />
                    <RANKING order="10" place="10" resultid="14134" />
                    <RANKING order="11" place="11" resultid="14422" />
                    <RANKING order="12" place="12" resultid="13967" />
                    <RANKING order="13" place="13" resultid="13377" />
                    <RANKING order="14" place="14" resultid="14273" />
                    <RANKING order="15" place="-1" resultid="14439" />
                    <RANKING order="16" place="-1" resultid="14344" />
                    <RANKING order="17" place="-1" resultid="12631" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14584" daytime="11:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14585" daytime="11:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14586" daytime="11:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14587" daytime="11:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14588" daytime="11:31" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14589" daytime="11:33" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1090" daytime="11:35" gender="M" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1147" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12774" />
                    <RANKING order="2" place="2" resultid="14158" />
                    <RANKING order="3" place="3" resultid="14083" />
                    <RANKING order="4" place="4" resultid="14127" />
                    <RANKING order="5" place="-1" resultid="14259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14030" />
                    <RANKING order="2" place="2" resultid="13032" />
                    <RANKING order="3" place="3" resultid="14512" />
                    <RANKING order="4" place="4" resultid="13329" />
                    <RANKING order="5" place="5" resultid="14404" />
                    <RANKING order="6" place="6" resultid="14070" />
                    <RANKING order="7" place="7" resultid="13325" />
                    <RANKING order="8" place="8" resultid="14337" />
                    <RANKING order="9" place="-1" resultid="14044" />
                    <RANKING order="10" place="-1" resultid="12694" />
                    <RANKING order="11" place="-1" resultid="13857" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14591" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14592" daytime="11:37" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14593" daytime="11:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14594" daytime="11:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="11:42" gender="F" number="13" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1164" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12783" />
                    <RANKING order="2" place="2" resultid="12135" />
                    <RANKING order="3" place="3" resultid="12707" />
                    <RANKING order="4" place="4" resultid="12119" />
                    <RANKING order="5" place="5" resultid="14025" />
                    <RANKING order="6" place="6" resultid="14340" />
                    <RANKING order="7" place="7" resultid="12914" />
                    <RANKING order="8" place="8" resultid="13319" />
                    <RANKING order="9" place="9" resultid="13014" />
                    <RANKING order="10" place="10" resultid="13148" />
                    <RANKING order="11" place="11" resultid="12502" />
                    <RANKING order="12" place="12" resultid="12788" />
                    <RANKING order="13" place="13" resultid="14351" />
                    <RANKING order="14" place="14" resultid="12801" />
                    <RANKING order="15" place="15" resultid="14215" />
                    <RANKING order="16" place="16" resultid="12749" />
                    <RANKING order="17" place="17" resultid="14062" />
                    <RANKING order="18" place="18" resultid="12115" />
                    <RANKING order="19" place="19" resultid="12805" />
                    <RANKING order="20" place="20" resultid="13809" />
                    <RANKING order="21" place="21" resultid="14393" />
                    <RANKING order="22" place="22" resultid="13916" />
                    <RANKING order="23" place="23" resultid="12489" />
                    <RANKING order="24" place="-1" resultid="12757" />
                    <RANKING order="25" place="-1" resultid="12900" />
                    <RANKING order="26" place="-1" resultid="13090" />
                    <RANKING order="27" place="-1" resultid="13267" />
                    <RANKING order="28" place="-1" resultid="13278" />
                    <RANKING order="29" place="-1" resultid="13875" />
                    <RANKING order="30" place="-1" resultid="13889" />
                    <RANKING order="31" place="-1" resultid="13920" />
                    <RANKING order="32" place="-1" resultid="14105" />
                    <RANKING order="33" place="-1" resultid="14373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13897" />
                    <RANKING order="2" place="2" resultid="12686" />
                    <RANKING order="3" place="3" resultid="12976" />
                    <RANKING order="4" place="4" resultid="13840" />
                    <RANKING order="5" place="5" resultid="13264" />
                    <RANKING order="6" place="6" resultid="12699" />
                    <RANKING order="7" place="7" resultid="13106" />
                    <RANKING order="8" place="8" resultid="13929" />
                    <RANKING order="9" place="9" resultid="14020" />
                    <RANKING order="10" place="10" resultid="12670" />
                    <RANKING order="11" place="11" resultid="12690" />
                    <RANKING order="12" place="12" resultid="12506" />
                    <RANKING order="13" place="13" resultid="14377" />
                    <RANKING order="14" place="14" resultid="12532" />
                    <RANKING order="15" place="15" resultid="12510" />
                    <RANKING order="16" place="16" resultid="13006" />
                    <RANKING order="17" place="17" resultid="13156" />
                    <RANKING order="18" place="-1" resultid="13027" />
                    <RANKING order="19" place="-1" resultid="13044" />
                    <RANKING order="20" place="-1" resultid="14246" />
                    <RANKING order="21" place="-1" resultid="12620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12892" />
                    <RANKING order="2" place="2" resultid="13196" />
                    <RANKING order="3" place="3" resultid="12921" />
                    <RANKING order="4" place="4" resultid="12933" />
                    <RANKING order="5" place="5" resultid="12815" />
                    <RANKING order="6" place="6" resultid="12745" />
                    <RANKING order="7" place="7" resultid="12704" />
                    <RANKING order="8" place="8" resultid="12547" />
                    <RANKING order="9" place="9" resultid="13296" />
                    <RANKING order="10" place="10" resultid="14431" />
                    <RANKING order="11" place="11" resultid="14035" />
                    <RANKING order="12" place="12" resultid="14242" />
                    <RANKING order="13" place="13" resultid="12963" />
                    <RANKING order="14" place="14" resultid="13193" />
                    <RANKING order="15" place="15" resultid="13056" />
                    <RANKING order="16" place="16" resultid="12575" />
                    <RANKING order="17" place="17" resultid="13833" />
                    <RANKING order="18" place="18" resultid="13972" />
                    <RANKING order="19" place="19" resultid="12178" />
                    <RANKING order="20" place="20" resultid="14362" />
                    <RANKING order="21" place="-1" resultid="14057" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14595" daytime="11:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14596" daytime="11:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14597" daytime="11:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14598" daytime="11:51" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14599" daytime="11:53" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14600" daytime="11:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14601" daytime="11:59" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14602" daytime="12:01" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14603" daytime="12:04" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14604" daytime="12:06" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14605" daytime="12:08" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14606" daytime="12:11" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14607" daytime="12:13" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14608" daytime="12:15" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14609" daytime="12:17" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14610" daytime="12:19" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="12:26" gender="M" number="14" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1167" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12793" />
                    <RANKING order="2" place="2" resultid="13076" />
                    <RANKING order="3" place="3" resultid="14053" />
                    <RANKING order="4" place="4" resultid="12570" />
                    <RANKING order="5" place="5" resultid="13257" />
                    <RANKING order="6" place="6" resultid="12753" />
                    <RANKING order="7" place="7" resultid="12537" />
                    <RANKING order="8" place="8" resultid="12761" />
                    <RANKING order="9" place="9" resultid="14100" />
                    <RANKING order="10" place="10" resultid="12718" />
                    <RANKING order="11" place="11" resultid="14180" />
                    <RANKING order="12" place="12" resultid="13805" />
                    <RANKING order="13" place="13" resultid="13048" />
                    <RANKING order="14" place="-1" resultid="12736" />
                    <RANKING order="15" place="-1" resultid="14114" />
                    <RANKING order="16" place="-1" resultid="14250" />
                    <RANKING order="17" place="-1" resultid="13136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12929" />
                    <RANKING order="2" place="2" resultid="14435" />
                    <RANKING order="3" place="3" resultid="12732" />
                    <RANKING order="4" place="4" resultid="14449" />
                    <RANKING order="5" place="5" resultid="13160" />
                    <RANKING order="6" place="6" resultid="13040" />
                    <RANKING order="7" place="7" resultid="13300" />
                    <RANKING order="8" place="8" resultid="14095" />
                    <RANKING order="9" place="9" resultid="12555" />
                    <RANKING order="10" place="10" resultid="12740" />
                    <RANKING order="11" place="11" resultid="14366" />
                    <RANKING order="12" place="12" resultid="13958" />
                    <RANKING order="13" place="13" resultid="13113" />
                    <RANKING order="14" place="14" resultid="12139" />
                    <RANKING order="15" place="15" resultid="12551" />
                    <RANKING order="16" place="16" resultid="14427" />
                    <RANKING order="17" place="17" resultid="12604" />
                    <RANKING order="18" place="18" resultid="14223" />
                    <RANKING order="19" place="-1" resultid="12797" />
                    <RANKING order="20" place="-1" resultid="13010" />
                    <RANKING order="21" place="-1" resultid="14118" />
                    <RANKING order="22" place="-1" resultid="13130" />
                    <RANKING order="23" place="-1" resultid="12612" />
                    <RANKING order="24" place="-1" resultid="13036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12714" />
                    <RANKING order="2" place="2" resultid="12968" />
                    <RANKING order="3" place="3" resultid="12904" />
                    <RANKING order="4" place="4" resultid="12810" />
                    <RANKING order="5" place="5" resultid="12864" />
                    <RANKING order="6" place="6" resultid="12728" />
                    <RANKING order="7" place="7" resultid="12896" />
                    <RANKING order="8" place="8" resultid="14166" />
                    <RANKING order="9" place="9" resultid="13316" />
                    <RANKING order="10" place="10" resultid="12170" />
                    <RANKING order="11" place="11" resultid="14171" />
                    <RANKING order="12" place="12" resultid="12770" />
                    <RANKING order="13" place="13" resultid="14066" />
                    <RANKING order="14" place="14" resultid="13954" />
                    <RANKING order="15" place="15" resultid="12639" />
                    <RANKING order="16" place="16" resultid="13816" />
                    <RANKING order="17" place="17" resultid="13370" />
                    <RANKING order="18" place="18" resultid="12765" />
                    <RANKING order="19" place="19" resultid="14154" />
                    <RANKING order="20" place="-1" resultid="12560" />
                    <RANKING order="21" place="-1" resultid="13052" />
                    <RANKING order="22" place="-1" resultid="13064" />
                    <RANKING order="23" place="-1" resultid="13366" />
                    <RANKING order="24" place="-1" resultid="13388" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14614" daytime="12:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14615" daytime="12:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14616" daytime="12:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14617" daytime="12:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14618" daytime="12:39" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14619" daytime="12:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14620" daytime="12:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14621" daytime="12:47" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14622" daytime="12:49" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14623" daytime="12:51" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14624" daytime="12:54" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14625" daytime="12:56" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14626" daytime="12:58" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14627" daytime="13:00" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14628" daytime="13:03" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14629" daytime="13:05" number="16" order="16" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1098" daytime="13:07" gender="F" number="15" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14822" />
                    <RANKING order="2" place="2" resultid="13872" />
                    <RANKING order="3" place="3" resultid="14017" />
                    <RANKING order="4" place="4" resultid="14397" />
                    <RANKING order="5" place="5" resultid="14228" />
                    <RANKING order="6" place="6" resultid="12609" />
                    <RANKING order="7" place="7" resultid="13913" />
                    <RANKING order="8" place="8" resultid="13854" />
                    <RANKING order="9" place="9" resultid="14151" />
                    <RANKING order="10" place="-1" resultid="12664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13020" />
                    <RANKING order="2" place="2" resultid="13082" />
                    <RANKING order="3" place="3" resultid="14124" />
                    <RANKING order="4" place="4" resultid="12724" />
                    <RANKING order="5" place="5" resultid="12960" />
                    <RANKING order="6" place="6" resultid="13902" />
                    <RANKING order="7" place="7" resultid="14238" />
                    <RANKING order="8" place="8" resultid="14386" />
                    <RANKING order="9" place="9" resultid="13968" />
                    <RANKING order="10" place="10" resultid="14423" />
                    <RANKING order="11" place="11" resultid="14135" />
                    <RANKING order="12" place="12" resultid="13378" />
                    <RANKING order="13" place="13" resultid="14440" />
                    <RANKING order="14" place="14" resultid="14049" />
                    <RANKING order="15" place="15" resultid="14002" />
                    <RANKING order="16" place="16" resultid="14274" />
                    <RANKING order="17" place="-1" resultid="14345" />
                    <RANKING order="18" place="-1" resultid="12632" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14631" daytime="13:07" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14632" daytime="13:09" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14633" daytime="13:11" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14634" daytime="13:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14635" daytime="13:13" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14636" daytime="13:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14637" daytime="13:16" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1100" daytime="13:18" gender="M" number="16" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1151" agemax="8" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14084" />
                    <RANKING order="2" place="2" resultid="12779" />
                    <RANKING order="3" place="3" resultid="12775" />
                    <RANKING order="4" place="4" resultid="14128" />
                    <RANKING order="5" place="5" resultid="14159" />
                    <RANKING order="6" place="-1" resultid="14260" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14031" />
                    <RANKING order="2" place="2" resultid="13033" />
                    <RANKING order="3" place="3" resultid="14510" />
                    <RANKING order="4" place="4" resultid="13328" />
                    <RANKING order="5" place="5" resultid="13326" />
                    <RANKING order="6" place="6" resultid="14405" />
                    <RANKING order="7" place="7" resultid="14336" />
                    <RANKING order="8" place="8" resultid="14045" />
                    <RANKING order="9" place="9" resultid="14071" />
                    <RANKING order="10" place="-1" resultid="12695" />
                    <RANKING order="11" place="-1" resultid="13858" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14638" daytime="13:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14639" daytime="13:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14640" daytime="13:21" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14641" daytime="13:22" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1102" daytime="13:25" gender="F" number="17" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1170" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14341" />
                    <RANKING order="2" place="2" resultid="12784" />
                    <RANKING order="3" place="3" resultid="12885" />
                    <RANKING order="4" place="4" resultid="12136" />
                    <RANKING order="5" place="5" resultid="12120" />
                    <RANKING order="6" place="6" resultid="14026" />
                    <RANKING order="7" place="7" resultid="14216" />
                    <RANKING order="8" place="8" resultid="13015" />
                    <RANKING order="9" place="9" resultid="12503" />
                    <RANKING order="10" place="10" resultid="12789" />
                    <RANKING order="11" place="11" resultid="14063" />
                    <RANKING order="12" place="12" resultid="14382" />
                    <RANKING order="13" place="13" resultid="13320" />
                    <RANKING order="14" place="14" resultid="12750" />
                    <RANKING order="15" place="15" resultid="12708" />
                    <RANKING order="16" place="16" resultid="12915" />
                    <RANKING order="17" place="17" resultid="13810" />
                    <RANKING order="18" place="18" resultid="13311" />
                    <RANKING order="19" place="18" resultid="14352" />
                    <RANKING order="20" place="20" resultid="13149" />
                    <RANKING order="21" place="21" resultid="12116" />
                    <RANKING order="22" place="22" resultid="12802" />
                    <RANKING order="23" place="23" resultid="13917" />
                    <RANKING order="24" place="24" resultid="14370" />
                    <RANKING order="25" place="25" resultid="14394" />
                    <RANKING order="26" place="26" resultid="12806" />
                    <RANKING order="27" place="27" resultid="14358" />
                    <RANKING order="28" place="28" resultid="12490" />
                    <RANKING order="29" place="-1" resultid="12758" />
                    <RANKING order="30" place="-1" resultid="12901" />
                    <RANKING order="31" place="-1" resultid="13091" />
                    <RANKING order="32" place="-1" resultid="13266" />
                    <RANKING order="33" place="-1" resultid="13279" />
                    <RANKING order="34" place="-1" resultid="13876" />
                    <RANKING order="35" place="-1" resultid="13890" />
                    <RANKING order="36" place="-1" resultid="13921" />
                    <RANKING order="37" place="-1" resultid="14106" />
                    <RANKING order="38" place="-1" resultid="14374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12687" />
                    <RANKING order="2" place="2" resultid="13841" />
                    <RANKING order="3" place="3" resultid="12691" />
                    <RANKING order="4" place="4" resultid="14378" />
                    <RANKING order="5" place="5" resultid="13898" />
                    <RANKING order="6" place="6" resultid="12700" />
                    <RANKING order="7" place="7" resultid="12977" />
                    <RANKING order="8" place="8" resultid="13930" />
                    <RANKING order="9" place="9" resultid="14021" />
                    <RANKING order="10" place="10" resultid="13045" />
                    <RANKING order="11" place="11" resultid="12533" />
                    <RANKING order="12" place="12" resultid="13307" />
                    <RANKING order="13" place="13" resultid="13007" />
                    <RANKING order="14" place="14" resultid="13107" />
                    <RANKING order="15" place="15" resultid="13157" />
                    <RANKING order="16" place="16" resultid="13263" />
                    <RANKING order="17" place="17" resultid="14247" />
                    <RANKING order="18" place="18" resultid="13294" />
                    <RANKING order="19" place="19" resultid="12507" />
                    <RANKING order="20" place="20" resultid="12511" />
                    <RANKING order="21" place="-1" resultid="13028" />
                    <RANKING order="22" place="-1" resultid="12148" />
                    <RANKING order="23" place="-1" resultid="12621" />
                    <RANKING order="24" place="-1" resultid="12671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12893" />
                    <RANKING order="2" place="2" resultid="14243" />
                    <RANKING order="3" place="3" resultid="13199" />
                    <RANKING order="4" place="4" resultid="12746" />
                    <RANKING order="5" place="5" resultid="12705" />
                    <RANKING order="6" place="6" resultid="14036" />
                    <RANKING order="7" place="7" resultid="12816" />
                    <RANKING order="8" place="8" resultid="12922" />
                    <RANKING order="9" place="9" resultid="12934" />
                    <RANKING order="10" place="10" resultid="13194" />
                    <RANKING order="11" place="11" resultid="12576" />
                    <RANKING order="12" place="12" resultid="12964" />
                    <RANKING order="13" place="13" resultid="13297" />
                    <RANKING order="14" place="14" resultid="13303" />
                    <RANKING order="15" place="15" resultid="13246" />
                    <RANKING order="16" place="16" resultid="12548" />
                    <RANKING order="17" place="16" resultid="13820" />
                    <RANKING order="18" place="18" resultid="13973" />
                    <RANKING order="19" place="19" resultid="14432" />
                    <RANKING order="20" place="20" resultid="13834" />
                    <RANKING order="21" place="21" resultid="13057" />
                    <RANKING order="22" place="22" resultid="14363" />
                    <RANKING order="23" place="23" resultid="12179" />
                    <RANKING order="24" place="24" resultid="13313" />
                    <RANKING order="25" place="-1" resultid="14058" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14643" daytime="13:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14644" daytime="13:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14645" daytime="13:31" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14646" daytime="13:33" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14647" daytime="13:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14648" daytime="13:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14649" daytime="13:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14650" daytime="13:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14651" daytime="13:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14652" daytime="13:46" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14653" daytime="13:48" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14654" daytime="13:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14655" daytime="13:52" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14656" daytime="13:54" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14657" daytime="13:56" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14658" daytime="13:57" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="14659" daytime="13:59" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="14660" daytime="14:01" number="18" order="18" status="OFFICIAL" />
                <HEAT heatid="14661" daytime="14:03" number="19" order="19" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="14:06" gender="M" number="18" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1174" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12930" />
                    <RANKING order="2" place="2" resultid="13161" />
                    <RANKING order="3" place="3" resultid="14119" />
                    <RANKING order="4" place="4" resultid="12733" />
                    <RANKING order="5" place="5" resultid="14450" />
                    <RANKING order="6" place="6" resultid="12798" />
                    <RANKING order="7" place="7" resultid="14367" />
                    <RANKING order="8" place="8" resultid="13299" />
                    <RANKING order="9" place="9" resultid="13959" />
                    <RANKING order="10" place="10" resultid="14224" />
                    <RANKING order="11" place="11" resultid="13011" />
                    <RANKING order="12" place="12" resultid="14096" />
                    <RANKING order="13" place="13" resultid="12741" />
                    <RANKING order="14" place="14" resultid="12140" />
                    <RANKING order="15" place="15" resultid="14436" />
                    <RANKING order="16" place="16" resultid="12556" />
                    <RANKING order="17" place="17" resultid="13041" />
                    <RANKING order="18" place="18" resultid="14428" />
                    <RANKING order="19" place="19" resultid="13131" />
                    <RANKING order="20" place="20" resultid="12613" />
                    <RANKING order="21" place="21" resultid="12605" />
                    <RANKING order="22" place="22" resultid="13114" />
                    <RANKING order="23" place="23" resultid="13910" />
                    <RANKING order="24" place="24" resultid="12552" />
                    <RANKING order="25" place="-1" resultid="13037" />
                    <RANKING order="26" place="-1" resultid="13285" />
                    <RANKING order="27" place="-1" resultid="13850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12794" />
                    <RANKING order="2" place="2" resultid="14101" />
                    <RANKING order="3" place="3" resultid="14054" />
                    <RANKING order="4" place="4" resultid="13077" />
                    <RANKING order="5" place="5" resultid="12719" />
                    <RANKING order="6" place="6" resultid="14181" />
                    <RANKING order="7" place="7" resultid="12571" />
                    <RANKING order="8" place="8" resultid="12754" />
                    <RANKING order="9" place="9" resultid="12538" />
                    <RANKING order="10" place="10" resultid="13806" />
                    <RANKING order="11" place="11" resultid="12737" />
                    <RANKING order="12" place="12" resultid="12762" />
                    <RANKING order="13" place="13" resultid="14115" />
                    <RANKING order="14" place="14" resultid="12911" />
                    <RANKING order="15" place="15" resultid="13049" />
                    <RANKING order="16" place="16" resultid="14251" />
                    <RANKING order="17" place="-1" resultid="13258" />
                    <RANKING order="18" place="-1" resultid="13946" />
                    <RANKING order="19" place="-1" resultid="13137" />
                    <RANKING order="20" place="-1" resultid="14401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12969" />
                    <RANKING order="2" place="2" resultid="14172" />
                    <RANKING order="3" place="3" resultid="12811" />
                    <RANKING order="4" place="4" resultid="12905" />
                    <RANKING order="5" place="5" resultid="13261" />
                    <RANKING order="6" place="6" resultid="12715" />
                    <RANKING order="7" place="7" resultid="12729" />
                    <RANKING order="8" place="8" resultid="12897" />
                    <RANKING order="9" place="9" resultid="12771" />
                    <RANKING order="10" place="10" resultid="12171" />
                    <RANKING order="11" place="11" resultid="14067" />
                    <RANKING order="12" place="12" resultid="13317" />
                    <RANKING order="13" place="13" resultid="13053" />
                    <RANKING order="14" place="14" resultid="13371" />
                    <RANKING order="15" place="15" resultid="12766" />
                    <RANKING order="16" place="16" resultid="13817" />
                    <RANKING order="17" place="17" resultid="12640" />
                    <RANKING order="18" place="18" resultid="12561" />
                    <RANKING order="19" place="19" resultid="13955" />
                    <RANKING order="20" place="20" resultid="14155" />
                    <RANKING order="21" place="-1" resultid="14167" />
                    <RANKING order="22" place="-1" resultid="12865" />
                    <RANKING order="23" place="-1" resultid="13943" />
                    <RANKING order="24" place="-1" resultid="13065" />
                    <RANKING order="25" place="-1" resultid="13367" />
                    <RANKING order="26" place="-1" resultid="13389" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14665" daytime="14:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14666" daytime="14:11" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14667" daytime="14:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14668" daytime="14:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14669" daytime="14:19" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14670" daytime="14:21" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14671" daytime="14:23" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14672" daytime="14:25" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14673" daytime="14:28" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14674" daytime="14:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14675" daytime="14:32" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14676" daytime="14:34" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14677" daytime="14:36" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14678" daytime="14:37" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14679" daytime="14:39" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14680" daytime="14:41" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="14681" daytime="14:43" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2022-12-03" daytime="16:30" endtime="17:58" name="De / Rü Nachmittag" number="5" warmupfrom="15:30" warmupuntil="16:20">
          <EVENTS>
            <EVENT eventid="1108" daytime="16:30" gender="F" number="21" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13084" />
                    <RANKING order="2" place="2" resultid="13163" />
                    <RANKING order="3" place="3" resultid="13937" />
                    <RANKING order="4" place="4" resultid="13254" />
                    <RANKING order="5" place="5" resultid="14230" />
                    <RANKING order="6" place="6" resultid="12181" />
                    <RANKING order="7" place="7" resultid="13093" />
                    <RANKING order="8" place="8" resultid="14354" />
                    <RANKING order="9" place="9" resultid="14446" />
                    <RANKING order="10" place="10" resultid="14412" />
                    <RANKING order="11" place="11" resultid="14108" />
                    <RANKING order="12" place="12" resultid="12521" />
                    <RANKING order="13" place="13" resultid="12492" />
                    <RANKING order="14" place="-1" resultid="12983" />
                    <RANKING order="15" place="-1" resultid="12859" />
                    <RANKING order="16" place="-1" resultid="12979" />
                    <RANKING order="17" place="-1" resultid="13181" />
                    <RANKING order="18" place="-1" resultid="13305" />
                    <RANKING order="19" place="-1" resultid="13383" />
                    <RANKING order="20" place="-1" resultid="14162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14004" />
                    <RANKING order="2" place="2" resultid="14077" />
                    <RANKING order="3" place="3" resultid="14038" />
                    <RANKING order="4" place="4" resultid="12879" />
                    <RANKING order="5" place="5" resultid="12871" />
                    <RANKING order="6" place="6" resultid="12186" />
                    <RANKING order="7" place="7" resultid="13865" />
                    <RANKING order="8" place="8" resultid="13187" />
                    <RANKING order="9" place="9" resultid="13290" />
                    <RANKING order="10" place="10" resultid="12154" />
                    <RANKING order="11" place="11" resultid="12526" />
                    <RANKING order="12" place="12" resultid="14140" />
                    <RANKING order="13" place="13" resultid="13883" />
                    <RANKING order="14" place="14" resultid="12517" />
                    <RANKING order="15" place="15" resultid="13116" />
                    <RANKING order="16" place="-1" resultid="12988" />
                    <RANKING order="17" place="-1" resultid="13948" />
                    <RANKING order="18" place="-1" resultid="14218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14267" />
                    <RANKING order="2" place="2" resultid="14276" />
                    <RANKING order="3" place="3" resultid="14193" />
                    <RANKING order="4" place="4" resultid="13961" />
                    <RANKING order="5" place="5" resultid="12165" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14684" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14685" daytime="16:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14686" daytime="16:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14687" daytime="16:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14688" daytime="16:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14689" daytime="16:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14690" daytime="16:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14691" daytime="16:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14692" daytime="16:45" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="16:49" gender="M" number="22" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1182" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14188" />
                    <RANKING order="2" place="2" resultid="14262" />
                    <RANKING order="3" place="3" resultid="14407" />
                    <RANKING order="4" place="4" resultid="12599" />
                    <RANKING order="5" place="5" resultid="14144" />
                    <RANKING order="6" place="6" resultid="13878" />
                    <RANKING order="7" place="7" resultid="13836" />
                    <RANKING order="8" place="8" resultid="12563" />
                    <RANKING order="9" place="-1" resultid="13373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13932" />
                    <RANKING order="2" place="2" resultid="12158" />
                    <RANKING order="3" place="3" resultid="14174" />
                    <RANKING order="4" place="4" resultid="13923" />
                    <RANKING order="5" place="5" resultid="14327" />
                    <RANKING order="6" place="6" resultid="14203" />
                    <RANKING order="7" place="7" resultid="12496" />
                    <RANKING order="8" place="-1" resultid="12992" />
                    <RANKING order="9" place="-1" resultid="13101" />
                    <RANKING order="10" place="-1" resultid="13391" />
                    <RANKING order="11" place="-1" resultid="14086" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14183" />
                    <RANKING order="2" place="2" resultid="13331" />
                    <RANKING order="3" place="3" resultid="13994" />
                    <RANKING order="4" place="4" resultid="13989" />
                    <RANKING order="5" place="5" resultid="14198" />
                    <RANKING order="6" place="6" resultid="12666" />
                    <RANKING order="7" place="7" resultid="13860" />
                    <RANKING order="8" place="8" resultid="14253" />
                    <RANKING order="9" place="9" resultid="13904" />
                    <RANKING order="10" place="10" resultid="12642" />
                    <RANKING order="11" place="-1" resultid="14208" />
                    <RANKING order="12" place="-1" resultid="14452" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14695" daytime="16:49" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14696" daytime="16:51" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14697" daytime="16:53" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14698" daytime="16:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14699" daytime="16:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14700" daytime="16:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14701" daytime="17:00" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="17:01" gender="F" number="23" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13086" />
                    <RANKING order="2" place="2" resultid="13938" />
                    <RANKING order="3" place="3" resultid="14109" />
                    <RANKING order="4" place="4" resultid="12142" />
                    <RANKING order="5" place="5" resultid="13164" />
                    <RANKING order="6" place="6" resultid="13178" />
                    <RANKING order="7" place="7" resultid="14355" />
                    <RANKING order="8" place="8" resultid="13022" />
                    <RANKING order="9" place="9" resultid="14137" />
                    <RANKING order="10" place="10" resultid="12182" />
                    <RANKING order="11" place="11" resultid="13094" />
                    <RANKING order="12" place="12" resultid="14231" />
                    <RANKING order="13" place="13" resultid="13201" />
                    <RANKING order="14" place="14" resultid="13001" />
                    <RANKING order="15" place="15" resultid="14012" />
                    <RANKING order="16" place="16" resultid="13287" />
                    <RANKING order="17" place="17" resultid="12522" />
                    <RANKING order="18" place="18" resultid="14413" />
                    <RANKING order="19" place="19" resultid="14443" />
                    <RANKING order="20" place="20" resultid="13812" />
                    <RANKING order="21" place="21" resultid="12650" />
                    <RANKING order="22" place="22" resultid="13269" />
                    <RANKING order="23" place="23" resultid="13126" />
                    <RANKING order="24" place="24" resultid="13122" />
                    <RANKING order="25" place="25" resultid="13151" />
                    <RANKING order="26" place="26" resultid="14417" />
                    <RANKING order="27" place="-1" resultid="13143" />
                    <RANKING order="28" place="-1" resultid="12984" />
                    <RANKING order="29" place="-1" resultid="13822" />
                    <RANKING order="30" place="-1" resultid="12860" />
                    <RANKING order="31" place="-1" resultid="12887" />
                    <RANKING order="32" place="-1" resultid="13380" />
                    <RANKING order="33" place="-1" resultid="13384" />
                    <RANKING order="34" place="-1" resultid="14073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13866" />
                    <RANKING order="2" place="2" resultid="14039" />
                    <RANKING order="3" place="3" resultid="14005" />
                    <RANKING order="4" place="4" resultid="14347" />
                    <RANKING order="5" place="5" resultid="14078" />
                    <RANKING order="6" place="6" resultid="12872" />
                    <RANKING order="7" place="7" resultid="13892" />
                    <RANKING order="8" place="8" resultid="12122" />
                    <RANKING order="9" place="9" resultid="12924" />
                    <RANKING order="10" place="10" resultid="14141" />
                    <RANKING order="11" place="11" resultid="12527" />
                    <RANKING order="12" place="12" resultid="12187" />
                    <RANKING order="13" place="13" resultid="12880" />
                    <RANKING order="14" place="14" resultid="13884" />
                    <RANKING order="15" place="15" resultid="13117" />
                    <RANKING order="16" place="16" resultid="14091" />
                    <RANKING order="17" place="17" resultid="12513" />
                    <RANKING order="18" place="-1" resultid="12658" />
                    <RANKING order="19" place="-1" resultid="12989" />
                    <RANKING order="20" place="-1" resultid="12634" />
                    <RANKING order="21" place="-1" resultid="13949" />
                    <RANKING order="22" place="-1" resultid="14219" />
                    <RANKING order="23" place="-1" resultid="14333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14268" />
                    <RANKING order="2" place="2" resultid="14194" />
                    <RANKING order="3" place="3" resultid="14277" />
                    <RANKING order="4" place="4" resultid="12166" />
                    <RANKING order="5" place="5" resultid="13962" />
                    <RANKING order="6" place="6" resultid="12126" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14703" daytime="17:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14704" daytime="17:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14705" daytime="17:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14706" daytime="17:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14707" daytime="17:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14708" daytime="17:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14709" daytime="17:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14710" daytime="17:15" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14711" daytime="17:17" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14712" daytime="17:19" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14713" daytime="17:21" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14714" daytime="17:22" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14715" daytime="17:24" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14716" daytime="17:26" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="17:29" gender="M" number="24" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1188" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14189" />
                    <RANKING order="2" place="2" resultid="13184" />
                    <RANKING order="3" place="3" resultid="14263" />
                    <RANKING order="4" place="4" resultid="13059" />
                    <RANKING order="5" place="5" resultid="12875" />
                    <RANKING order="6" place="6" resultid="14408" />
                    <RANKING order="7" place="7" resultid="12867" />
                    <RANKING order="8" place="8" resultid="13098" />
                    <RANKING order="9" place="9" resultid="14145" />
                    <RANKING order="10" place="10" resultid="13139" />
                    <RANKING order="11" place="11" resultid="13879" />
                    <RANKING order="12" place="12" resultid="12615" />
                    <RANKING order="13" place="13" resultid="12150" />
                    <RANKING order="14" place="14" resultid="12971" />
                    <RANKING order="15" place="15" resultid="12564" />
                    <RANKING order="16" place="16" resultid="12173" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12159" />
                    <RANKING order="2" place="2" resultid="13933" />
                    <RANKING order="3" place="3" resultid="14328" />
                    <RANKING order="4" place="4" resultid="12646" />
                    <RANKING order="5" place="5" resultid="13924" />
                    <RANKING order="6" place="6" resultid="12917" />
                    <RANKING order="7" place="7" resultid="14204" />
                    <RANKING order="8" place="8" resultid="14175" />
                    <RANKING order="9" place="9" resultid="12997" />
                    <RANKING order="10" place="10" resultid="12907" />
                    <RANKING order="11" place="11" resultid="12654" />
                    <RANKING order="12" place="12" resultid="13251" />
                    <RANKING order="13" place="13" resultid="12623" />
                    <RANKING order="14" place="-1" resultid="12130" />
                    <RANKING order="15" place="-1" resultid="12993" />
                    <RANKING order="16" place="-1" resultid="13070" />
                    <RANKING order="17" place="-1" resultid="13102" />
                    <RANKING order="18" place="-1" resultid="14087" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14184" />
                    <RANKING order="2" place="2" resultid="13995" />
                    <RANKING order="3" place="3" resultid="14199" />
                    <RANKING order="4" place="4" resultid="14453" />
                    <RANKING order="5" place="5" resultid="13861" />
                    <RANKING order="6" place="6" resultid="13905" />
                    <RANKING order="7" place="7" resultid="14254" />
                    <RANKING order="8" place="8" resultid="12643" />
                    <RANKING order="9" place="9" resultid="13990" />
                    <RANKING order="10" place="-1" resultid="13322" />
                    <RANKING order="11" place="-1" resultid="14130" />
                    <RANKING order="12" place="-1" resultid="14209" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14719" daytime="17:29" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14720" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14721" daytime="17:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14722" daytime="17:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14723" daytime="17:37" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14724" daytime="17:39" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14725" daytime="17:41" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14726" daytime="17:43" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14727" daytime="17:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14728" daytime="17:46" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14729" daytime="17:47" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2022-12-03" daytime="17:56" endtime="18:11" name="Staffeln Lagen Nachmittag" number="6">
          <EVENTS>
            <EVENT eventid="1120" daytime="17:56" gender="F" number="25" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="CHF" value="1800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1121" agemax="-1" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14285" />
                    <RANKING order="2" place="2" resultid="12189" />
                    <RANKING order="3" place="3" resultid="13976" />
                    <RANKING order="4" place="4" resultid="14458" />
                    <RANKING order="5" place="5" resultid="13172" />
                    <RANKING order="6" place="6" resultid="14287" />
                    <RANKING order="7" place="7" resultid="13174" />
                    <RANKING order="8" place="8" resultid="12579" />
                    <RANKING order="9" place="9" resultid="13336" />
                    <RANKING order="10" place="-1" resultid="14286" />
                    <RANKING order="11" place="-1" resultid="12938" />
                    <RANKING order="12" place="-1" resultid="13203" />
                    <RANKING order="13" place="-1" resultid="13338" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14731" daytime="17:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14732" daytime="17:59" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14733" daytime="18:02" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="18:05" gender="M" number="26" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="CHF" value="1800" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="-1" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14283" />
                    <RANKING order="2" place="2" resultid="13975" />
                    <RANKING order="3" place="3" resultid="12672" />
                    <RANKING order="4" place="4" resultid="14284" />
                    <RANKING order="5" place="5" resultid="13334" />
                    <RANKING order="6" place="6" resultid="13168" />
                    <RANKING order="7" place="7" resultid="12936" />
                    <RANKING order="8" place="8" resultid="12673" />
                    <RANKING order="9" place="-1" resultid="13170" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14735" daytime="18:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14736" daytime="18:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2022-12-03" daytime="18:18" endtime="19:53" name="Br / Cr Nachmittag" number="7">
          <EVENTS>
            <EVENT eventid="1124" daytime="18:18" gender="F" number="27" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1191" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12143" />
                    <RANKING order="2" place="2" resultid="13939" />
                    <RANKING order="3" place="3" resultid="14444" />
                    <RANKING order="4" place="4" resultid="13002" />
                    <RANKING order="5" place="5" resultid="14389" />
                    <RANKING order="6" place="6" resultid="14110" />
                    <RANKING order="7" place="7" resultid="13095" />
                    <RANKING order="8" place="8" resultid="12183" />
                    <RANKING order="9" place="9" resultid="13085" />
                    <RANKING order="10" place="10" resultid="13273" />
                    <RANKING order="11" place="11" resultid="13144" />
                    <RANKING order="12" place="12" resultid="14013" />
                    <RANKING order="13" place="13" resultid="13023" />
                    <RANKING order="14" place="14" resultid="13275" />
                    <RANKING order="15" place="15" resultid="12523" />
                    <RANKING order="16" place="16" resultid="12493" />
                    <RANKING order="17" place="17" resultid="12651" />
                    <RANKING order="18" place="18" resultid="13152" />
                    <RANKING order="19" place="19" resultid="14414" />
                    <RANKING order="20" place="20" resultid="13127" />
                    <RANKING order="21" place="21" resultid="13123" />
                    <RANKING order="22" place="22" resultid="14418" />
                    <RANKING order="23" place="-1" resultid="13165" />
                    <RANKING order="24" place="-1" resultid="12985" />
                    <RANKING order="25" place="-1" resultid="12888" />
                    <RANKING order="26" place="-1" resultid="12980" />
                    <RANKING order="27" place="-1" resultid="14074" />
                    <RANKING order="28" place="-1" resultid="14232" />
                    <RANKING order="29" place="-1" resultid="14161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14079" />
                    <RANKING order="2" place="2" resultid="13983" />
                    <RANKING order="3" place="3" resultid="14006" />
                    <RANKING order="4" place="4" resultid="12155" />
                    <RANKING order="5" place="5" resultid="14281" />
                    <RANKING order="6" place="6" resultid="14040" />
                    <RANKING order="7" place="7" resultid="13867" />
                    <RANKING order="8" place="8" resultid="12123" />
                    <RANKING order="9" place="9" resultid="12518" />
                    <RANKING order="10" place="10" resultid="13893" />
                    <RANKING order="11" place="11" resultid="13885" />
                    <RANKING order="12" place="12" resultid="12925" />
                    <RANKING order="13" place="13" resultid="14092" />
                    <RANKING order="14" place="14" resultid="13281" />
                    <RANKING order="15" place="15" resultid="12528" />
                    <RANKING order="16" place="16" resultid="13109" />
                    <RANKING order="17" place="17" resultid="12514" />
                    <RANKING order="18" place="18" resultid="12659" />
                    <RANKING order="19" place="19" resultid="12162" />
                    <RANKING order="20" place="-1" resultid="13118" />
                    <RANKING order="21" place="-1" resultid="12635" />
                    <RANKING order="22" place="-1" resultid="13950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14269" />
                    <RANKING order="2" place="2" resultid="14009" />
                    <RANKING order="3" place="3" resultid="14278" />
                    <RANKING order="4" place="4" resultid="14195" />
                    <RANKING order="5" place="5" resultid="13963" />
                    <RANKING order="6" place="6" resultid="12127" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14738" daytime="18:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14739" daytime="18:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14740" daytime="18:23" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14741" daytime="18:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14742" daytime="18:27" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14743" daytime="18:29" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14744" daytime="18:31" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14745" daytime="18:33" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14746" daytime="18:35" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14747" daytime="18:37" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14748" daytime="18:39" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14749" daytime="18:41" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14750" daytime="18:43" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" daytime="18:47" gender="M" number="28" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1194" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14190" />
                    <RANKING order="2" place="2" resultid="14409" />
                    <RANKING order="3" place="3" resultid="14264" />
                    <RANKING order="4" place="4" resultid="12876" />
                    <RANKING order="5" place="5" resultid="12868" />
                    <RANKING order="6" place="6" resultid="13060" />
                    <RANKING order="7" place="7" resultid="13140" />
                    <RANKING order="8" place="8" resultid="12600" />
                    <RANKING order="9" place="9" resultid="12616" />
                    <RANKING order="10" place="10" resultid="13880" />
                    <RANKING order="11" place="11" resultid="12151" />
                    <RANKING order="12" place="12" resultid="12174" />
                    <RANKING order="13" place="13" resultid="12972" />
                    <RANKING order="14" place="14" resultid="12565" />
                    <RANKING order="15" place="-1" resultid="14146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13986" />
                    <RANKING order="2" place="2" resultid="13925" />
                    <RANKING order="3" place="3" resultid="13934" />
                    <RANKING order="4" place="4" resultid="13248" />
                    <RANKING order="5" place="5" resultid="12647" />
                    <RANKING order="6" place="6" resultid="13190" />
                    <RANKING order="7" place="7" resultid="14329" />
                    <RANKING order="8" place="8" resultid="14205" />
                    <RANKING order="9" place="9" resultid="14176" />
                    <RANKING order="10" place="10" resultid="13067" />
                    <RANKING order="11" place="11" resultid="12497" />
                    <RANKING order="12" place="12" resultid="12998" />
                    <RANKING order="13" place="13" resultid="12624" />
                    <RANKING order="14" place="14" resultid="13825" />
                    <RANKING order="15" place="15" resultid="12131" />
                    <RANKING order="16" place="-1" resultid="12655" />
                    <RANKING order="17" place="-1" resultid="12994" />
                    <RANKING order="18" place="-1" resultid="13071" />
                    <RANKING order="19" place="-1" resultid="14088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12856" />
                    <RANKING order="2" place="2" resultid="13996" />
                    <RANKING order="3" place="3" resultid="14200" />
                    <RANKING order="4" place="4" resultid="14185" />
                    <RANKING order="5" place="5" resultid="12627" />
                    <RANKING order="6" place="6" resultid="13991" />
                    <RANKING order="7" place="7" resultid="13906" />
                    <RANKING order="8" place="8" resultid="13862" />
                    <RANKING order="9" place="9" resultid="14255" />
                    <RANKING order="10" place="-1" resultid="14131" />
                    <RANKING order="11" place="-1" resultid="14210" />
                    <RANKING order="12" place="-1" resultid="14454" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14753" daytime="18:47" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14754" daytime="18:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14755" daytime="18:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14756" daytime="18:53" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14757" daytime="18:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14758" daytime="18:57" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14759" daytime="18:59" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14760" daytime="19:01" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14761" daytime="19:03" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14762" daytime="19:04" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14763" daytime="19:06" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="19:08" gender="F" number="29" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13087" />
                    <RANKING order="2" place="2" resultid="13940" />
                    <RANKING order="3" place="3" resultid="12144" />
                    <RANKING order="4" place="4" resultid="13179" />
                    <RANKING order="5" place="5" resultid="14111" />
                    <RANKING order="6" place="6" resultid="14390" />
                    <RANKING order="7" place="7" resultid="14356" />
                    <RANKING order="8" place="8" resultid="12184" />
                    <RANKING order="9" place="9" resultid="14233" />
                    <RANKING order="10" place="10" resultid="14138" />
                    <RANKING order="11" place="11" resultid="13166" />
                    <RANKING order="12" place="12" resultid="13255" />
                    <RANKING order="13" place="13" resultid="13096" />
                    <RANKING order="14" place="14" resultid="14445" />
                    <RANKING order="15" place="15" resultid="13024" />
                    <RANKING order="16" place="16" resultid="13003" />
                    <RANKING order="17" place="17" resultid="13145" />
                    <RANKING order="18" place="18" resultid="14415" />
                    <RANKING order="19" place="19" resultid="13276" />
                    <RANKING order="20" place="20" resultid="13270" />
                    <RANKING order="21" place="21" resultid="12652" />
                    <RANKING order="22" place="22" resultid="12524" />
                    <RANKING order="23" place="23" resultid="13288" />
                    <RANKING order="24" place="24" resultid="13202" />
                    <RANKING order="25" place="25" resultid="13813" />
                    <RANKING order="26" place="26" resultid="12494" />
                    <RANKING order="27" place="27" resultid="13124" />
                    <RANKING order="28" place="28" resultid="13128" />
                    <RANKING order="29" place="29" resultid="14419" />
                    <RANKING order="30" place="30" resultid="13153" />
                    <RANKING order="31" place="-1" resultid="12986" />
                    <RANKING order="32" place="-1" resultid="13823" />
                    <RANKING order="33" place="-1" resultid="12861" />
                    <RANKING order="34" place="-1" resultid="12889" />
                    <RANKING order="35" place="-1" resultid="12981" />
                    <RANKING order="36" place="-1" resultid="13182" />
                    <RANKING order="37" place="-1" resultid="13381" />
                    <RANKING order="38" place="-1" resultid="13385" />
                    <RANKING order="39" place="-1" resultid="14075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14007" />
                    <RANKING order="2" place="2" resultid="14080" />
                    <RANKING order="3" place="3" resultid="13868" />
                    <RANKING order="4" place="4" resultid="12124" />
                    <RANKING order="5" place="5" resultid="13984" />
                    <RANKING order="6" place="6" resultid="12188" />
                    <RANKING order="7" place="6" resultid="14041" />
                    <RANKING order="8" place="8" resultid="13894" />
                    <RANKING order="9" place="9" resultid="14348" />
                    <RANKING order="10" place="10" resultid="12881" />
                    <RANKING order="11" place="11" resultid="12873" />
                    <RANKING order="12" place="12" resultid="13188" />
                    <RANKING order="13" place="13" resultid="12529" />
                    <RANKING order="14" place="14" resultid="12156" />
                    <RANKING order="15" place="15" resultid="14282" />
                    <RANKING order="16" place="16" resultid="13291" />
                    <RANKING order="17" place="17" resultid="14142" />
                    <RANKING order="18" place="18" resultid="13886" />
                    <RANKING order="19" place="19" resultid="12519" />
                    <RANKING order="20" place="20" resultid="13119" />
                    <RANKING order="21" place="21" resultid="12926" />
                    <RANKING order="22" place="22" resultid="13282" />
                    <RANKING order="23" place="23" resultid="13110" />
                    <RANKING order="24" place="24" resultid="12163" />
                    <RANKING order="25" place="25" resultid="12660" />
                    <RANKING order="26" place="26" resultid="12515" />
                    <RANKING order="27" place="-1" resultid="12990" />
                    <RANKING order="28" place="-1" resultid="12636" />
                    <RANKING order="29" place="-1" resultid="13951" />
                    <RANKING order="30" place="-1" resultid="14220" />
                    <RANKING order="31" place="-1" resultid="14332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14270" />
                    <RANKING order="2" place="2" resultid="14279" />
                    <RANKING order="3" place="3" resultid="14196" />
                    <RANKING order="4" place="4" resultid="14288" />
                    <RANKING order="5" place="5" resultid="12167" />
                    <RANKING order="6" place="6" resultid="13964" />
                    <RANKING order="7" place="7" resultid="12128" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14765" daytime="19:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14766" daytime="19:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14767" daytime="19:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14768" daytime="19:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14769" daytime="19:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14770" daytime="19:17" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14771" daytime="19:19" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14772" daytime="19:21" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14773" daytime="19:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14774" daytime="19:24" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14775" daytime="19:26" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14776" daytime="19:27" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14777" daytime="19:29" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14778" daytime="19:30" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="14779" daytime="19:32" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="14780" daytime="19:33" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="14781" daytime="19:35" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1133" daytime="19:38" gender="M" number="30" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1199" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13987" />
                    <RANKING order="2" place="2" resultid="12160" />
                    <RANKING order="3" place="3" resultid="13935" />
                    <RANKING order="4" place="4" resultid="12918" />
                    <RANKING order="5" place="5" resultid="13926" />
                    <RANKING order="6" place="6" resultid="14177" />
                    <RANKING order="7" place="7" resultid="13191" />
                    <RANKING order="8" place="8" resultid="14206" />
                    <RANKING order="9" place="9" resultid="12648" />
                    <RANKING order="10" place="10" resultid="14330" />
                    <RANKING order="11" place="11" resultid="12625" />
                    <RANKING order="12" place="12" resultid="12498" />
                    <RANKING order="13" place="13" resultid="13252" />
                    <RANKING order="14" place="14" resultid="13068" />
                    <RANKING order="15" place="15" resultid="12999" />
                    <RANKING order="16" place="16" resultid="12908" />
                    <RANKING order="17" place="17" resultid="13249" />
                    <RANKING order="18" place="18" resultid="12656" />
                    <RANKING order="19" place="19" resultid="13826" />
                    <RANKING order="20" place="20" resultid="12132" />
                    <RANKING order="21" place="-1" resultid="12995" />
                    <RANKING order="22" place="-1" resultid="13072" />
                    <RANKING order="23" place="-1" resultid="13103" />
                    <RANKING order="24" place="-1" resultid="13392" />
                    <RANKING order="25" place="-1" resultid="14089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14191" />
                    <RANKING order="2" place="2" resultid="14265" />
                    <RANKING order="3" place="3" resultid="13185" />
                    <RANKING order="4" place="4" resultid="14410" />
                    <RANKING order="5" place="5" resultid="12877" />
                    <RANKING order="6" place="6" resultid="12869" />
                    <RANKING order="7" place="7" resultid="13061" />
                    <RANKING order="8" place="8" resultid="13099" />
                    <RANKING order="9" place="9" resultid="12601" />
                    <RANKING order="10" place="10" resultid="14147" />
                    <RANKING order="11" place="11" resultid="12152" />
                    <RANKING order="12" place="12" resultid="12617" />
                    <RANKING order="13" place="13" resultid="13141" />
                    <RANKING order="14" place="14" resultid="13837" />
                    <RANKING order="15" place="15" resultid="13881" />
                    <RANKING order="16" place="16" resultid="12973" />
                    <RANKING order="17" place="17" resultid="12175" />
                    <RANKING order="18" place="18" resultid="12566" />
                    <RANKING order="19" place="-1" resultid="13374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14455" />
                    <RANKING order="2" place="2" resultid="14186" />
                    <RANKING order="3" place="3" resultid="12854" />
                    <RANKING order="4" place="4" resultid="13997" />
                    <RANKING order="5" place="5" resultid="13332" />
                    <RANKING order="6" place="6" resultid="14201" />
                    <RANKING order="7" place="7" resultid="13992" />
                    <RANKING order="8" place="8" resultid="12667" />
                    <RANKING order="9" place="9" resultid="12644" />
                    <RANKING order="10" place="10" resultid="13863" />
                    <RANKING order="11" place="11" resultid="14256" />
                    <RANKING order="12" place="12" resultid="13907" />
                    <RANKING order="13" place="13" resultid="12628" />
                    <RANKING order="14" place="14" resultid="13323" />
                    <RANKING order="15" place="-1" resultid="14211" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14784" daytime="19:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14785" daytime="19:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14786" daytime="19:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14787" daytime="19:43" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14788" daytime="19:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="14789" daytime="19:47" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14790" daytime="19:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14791" daytime="19:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14792" daytime="19:51" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="14793" daytime="19:53" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="14794" daytime="19:54" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="14795" daytime="19:55" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="14796" daytime="19:57" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="14797" daytime="19:58" number="14" order="14" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2022-12-03" daytime="20:10" name="Sprint Cup" number="8">
          <EVENTS>
            <EVENT eventid="6685" daytime="20:10" gender="F" number="101" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6686" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14845" />
                    <RANKING order="2" place="2" resultid="14846" />
                    <RANKING order="3" place="3" resultid="14844" />
                    <RANKING order="4" place="4" resultid="14849" />
                    <RANKING order="5" place="5" resultid="14850" />
                    <RANKING order="6" place="6" resultid="14847" />
                    <RANKING order="7" place="7" resultid="14851" />
                    <RANKING order="8" place="8" resultid="14848" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14801" daytime="20:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14842" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6687" daytime="20:14" gender="M" number="102" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6688" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14854" />
                    <RANKING order="2" place="2" resultid="14858" />
                    <RANKING order="3" place="3" resultid="14857" />
                    <RANKING order="4" place="4" resultid="14859" />
                    <RANKING order="5" place="5" resultid="14856" />
                    <RANKING order="6" place="6" resultid="14852" />
                    <RANKING order="7" place="7" resultid="14855" />
                    <RANKING order="8" place="8" resultid="14853" />
                    <RANKING order="9" place="-1" resultid="14495" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14802" daytime="20:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14843" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14861" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6681" daytime="20:17" gender="F" number="103" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6682" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14862" />
                    <RANKING order="2" place="2" resultid="14864" />
                    <RANKING order="3" place="3" resultid="14863" />
                    <RANKING order="4" place="4" resultid="14865" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14803" daytime="20:17" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6683" daytime="20:21" gender="M" number="104" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6684" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14866" />
                    <RANKING order="2" place="2" resultid="14869" />
                    <RANKING order="3" place="3" resultid="14868" />
                    <RANKING order="4" place="4" resultid="14867" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14804" daytime="20:21" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6635" daytime="20:24" gender="F" number="105" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6636" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14870" />
                    <RANKING order="2" place="2" resultid="14871" />
                    <RANKING order="3" place="3" resultid="14872" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14805" daytime="20:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6639" daytime="20:28" gender="M" number="106" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6640" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14873" />
                    <RANKING order="2" place="2" resultid="14875" />
                    <RANKING order="3" place="3" resultid="14874" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14806" daytime="20:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6637" daytime="20:31" gender="F" number="107" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6638" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14876" />
                    <RANKING order="2" place="2" resultid="14877" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14807" daytime="20:31" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="6679" daytime="20:35" gender="M" number="108" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6680" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14878" />
                    <RANKING order="2" place="2" resultid="14879" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="14808" daytime="20:35" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14834" role="REF" />
          </JUDGES>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="SRM" nation="SUI" region="RSR" clubid="12112" swrid="65709" name="Schwimmklub Region Murten" shortname="Srm">
          <ATHLETES>
            <ATHLETE firstname="Janina" lastname="Zürcher" birthdate="2009-05-01" gender="F" nation="SUI" license="3618" swrid="4415945" athleteid="12180">
              <RESULTS>
                <RESULT eventid="1108" points="281" swimtime="00:01:23.37" resultid="12181" heatid="14687" lane="4" entrytime="00:01:28.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="75" swimtime="00:00:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="308" swimtime="00:01:21.23" resultid="12182" heatid="14710" lane="1" entrytime="00:01:20.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.72" />
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="75" swimtime="00:01:01.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="321" swimtime="00:01:31.04" resultid="12183" heatid="14745" lane="1" entrytime="00:01:30.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.50" />
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                    <SPLIT distance="75" swimtime="00:01:07.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="392" swimtime="00:01:08.65" resultid="12184" heatid="14774" lane="3" entrytime="00:01:08.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.58" />
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="75" swimtime="00:00:51.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maximilien" lastname="Salathé" birthdate="2008-09-05" gender="M" nation="SUI" license="42282" swrid="5559294" athleteid="12172">
              <RESULTS>
                <RESULT eventid="1117" points="107" swimtime="00:01:41.51" resultid="12173" heatid="14719" lane="1" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.61" />
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="75" swimtime="00:01:14.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="149" swimtime="00:01:44.34" resultid="12174" heatid="14753" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.53" />
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                    <SPLIT distance="75" swimtime="00:01:15.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="147" swimtime="00:01:24.97" resultid="12175" heatid="14784" lane="2" entrytime="00:01:24.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.14" />
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luc" lastname="Mathys" birthdate="2006-11-17" gender="M" nation="SUI" license="3627" swrid="5297935" athleteid="12157">
              <RESULTS>
                <RESULT eventid="1111" points="419" swimtime="00:01:03.81" resultid="12158" heatid="14700" lane="4" entrytime="00:01:04.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.07" />
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="75" swimtime="00:00:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="356" swimtime="00:01:08.13" resultid="12159" heatid="14728" lane="4" entrytime="00:01:07.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:50.70" />
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="528" swimtime="00:00:55.57" resultid="12160" heatid="14796" lane="1" entrytime="00:00:55.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.53" />
                    <SPLIT distance="50" swimtime="00:00:26.20" />
                    <SPLIT distance="75" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="369" swimtime="00:00:30.96" resultid="14855" heatid="14802" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nives" lastname="Blatter" birthdate="2011-07-31" gender="F" nation="SUI" license="32532" swrid="5466254" athleteid="12117">
              <RESULTS>
                <RESULT eventid="1078" points="246" swimtime="00:01:27.50" resultid="12118" heatid="14552" lane="4" entrytime="00:01:33.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.01" />
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="272" swimtime="00:01:36.20" resultid="12119" heatid="14607" lane="1" entrytime="00:01:41.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.79" />
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                    <SPLIT distance="75" swimtime="00:01:11.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="286" swimtime="00:01:16.19" resultid="12120" heatid="14658" lane="2" entrytime="00:01:17.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.66" />
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="75" swimtime="00:00:57.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malin" lastname="Kocher" birthdate="2012-02-19" gender="F" nation="SUI" license="3630" swrid="4403611" athleteid="12145">
              <RESULTS>
                <RESULT eventid="1068" status="WDR" swimtime="00:00:00.00" resultid="12146" entrytime="00:01:34.47" entrycourse="SCM" />
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="12147" entrytime="00:01:33.42" entrycourse="LCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="12148" entrytime="00:01:13.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Loïc" lastname="Hersberger" birthdate="2012-12-29" gender="M" nation="SUI" license="42280" swrid="5559911" athleteid="12137">
              <RESULTS>
                <RESULT eventid="1081" points="63" swimtime="00:02:01.42" resultid="12138" heatid="14567" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.70" />
                    <SPLIT distance="50" swimtime="00:00:58.41" />
                    <SPLIT distance="75" swimtime="00:01:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="72" swimtime="00:02:13.01" resultid="12139" heatid="14623" lane="3" entrytime="00:01:53.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.60" />
                    <SPLIT distance="50" swimtime="00:01:02.34" />
                    <SPLIT distance="75" swimtime="00:01:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="91" swimtime="00:01:39.72" resultid="12140" heatid="14670" lane="2" entrytime="00:01:41.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.38" />
                    <SPLIT distance="50" swimtime="00:00:45.81" />
                    <SPLIT distance="75" swimtime="00:01:14.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Louis" lastname="Herren" birthdate="2007-12-30" gender="M" nation="SUI" license="42284" swrid="5559290" athleteid="12129">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 17:39)" eventid="1117" status="DSQ" swimtime="00:01:40.31" resultid="12130" heatid="14719" lane="3" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.98" />
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="170" swimtime="00:01:39.79" resultid="12131" heatid="14753" lane="2" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.05" />
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                    <SPLIT distance="75" swimtime="00:01:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="202" swimtime="00:01:16.47" resultid="12132" heatid="14784" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.22" />
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="75" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livio" lastname="Reusser" birthdate="2010-05-28" gender="M" nation="SUI" license="42283" swrid="5559292" athleteid="12168">
              <RESULTS>
                <RESULT eventid="1081" points="117" swimtime="00:01:38.56" resultid="12169" heatid="14568" lane="3" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.29" />
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                    <SPLIT distance="75" swimtime="00:01:14.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="144" swimtime="00:01:45.56" resultid="12170" heatid="14624" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.82" />
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                    <SPLIT distance="75" swimtime="00:01:19.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="134" swimtime="00:01:27.66" resultid="12171" heatid="14675" lane="4" entrytime="00:01:32.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.34" />
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                    <SPLIT distance="75" swimtime="00:01:06.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noemi Anna" lastname="Marti" birthdate="2007-03-02" gender="F" nation="SUI" license="3635" swrid="5297918" athleteid="12153">
              <RESULTS>
                <RESULT eventid="1108" points="297" swimtime="00:01:21.79" resultid="12154" heatid="14687" lane="3" entrytime="00:01:25.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.46" />
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="75" swimtime="00:00:57.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="430" swimtime="00:01:22.58" resultid="12155" heatid="14747" lane="2" entrytime="00:01:24.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.32" />
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="75" swimtime="00:01:00.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="396" swimtime="00:01:08.38" resultid="12156" heatid="14776" lane="1" entrytime="00:01:06.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.22" />
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="75" swimtime="00:00:50.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Morgane" lastname="Degoumois" birthdate="2005-09-10" gender="F" nation="SUI" license="3632" swrid="5326602" athleteid="12125">
              <RESULTS>
                <RESULT eventid="1114" points="281" swimtime="00:01:23.76" resultid="12126" heatid="14706" lane="2" entrytime="00:01:29.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.61" />
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="261" swimtime="00:01:37.46" resultid="12127" heatid="14740" lane="2" entrytime="00:01:41.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.42" />
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                    <SPLIT distance="75" swimtime="00:01:11.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="355" swimtime="00:01:10.92" resultid="12128" heatid="14772" lane="3" entrytime="00:01:11.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.47" />
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="75" swimtime="00:00:53.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Josephine" lastname="Ober" birthdate="2007-04-29" gender="F" nation="SUI" license="42289" swrid="5559291" athleteid="12161">
              <RESULTS>
                <RESULT eventid="1124" points="153" swimtime="00:01:56.35" resultid="12162" heatid="14738" lane="2" entrytime="00:01:56.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.67" />
                    <SPLIT distance="50" swimtime="00:00:52.94" />
                    <SPLIT distance="75" swimtime="00:01:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="200" swimtime="00:01:25.81" resultid="12163" heatid="14766" lane="3" entrytime="00:01:28.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.86" />
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="75" swimtime="00:01:03.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leoni" lastname="Petersen" birthdate="2004-12-09" gender="F" nation="GER" license="3624" swrid="4971866" athleteid="12164">
              <RESULTS>
                <RESULT eventid="1108" points="321" swimtime="00:01:19.71" resultid="12165" heatid="14688" lane="4" entrytime="00:01:23.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="75" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="344" swimtime="00:01:18.27" resultid="12166" heatid="14712" lane="2" entrytime="00:01:17.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.44" />
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                    <SPLIT distance="75" swimtime="00:00:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="459" swimtime="00:01:05.14" resultid="12167" heatid="14778" lane="2" entrytime="00:01:04.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.66" />
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="75" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphaël" lastname="Marcolino" birthdate="2008-08-19" gender="M" nation="SUI" license="34880" swrid="5168734" athleteid="12149">
              <RESULTS>
                <RESULT eventid="1117" points="152" swimtime="00:01:30.45" resultid="12150" heatid="14720" lane="2" entrytime="00:01:29.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="174" swimtime="00:01:39.08" resultid="12151" heatid="14754" lane="2" entrytime="00:01:44.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.50" />
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="75" swimtime="00:01:11.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="243" swimtime="00:01:12.00" resultid="12152" heatid="14785" lane="3" entrytime="00:01:16.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.60" />
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="75" swimtime="00:00:53.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leah" lastname="Kocher" birthdate="2009-12-24" gender="F" nation="SUI" license="3623" swrid="4568526" athleteid="12141">
              <RESULTS>
                <RESULT eventid="1114" points="360" swimtime="00:01:17.12" resultid="12142" heatid="14711" lane="2" entrytime="00:01:18.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.10" />
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                    <SPLIT distance="75" swimtime="00:00:57.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="475" swimtime="00:01:19.90" resultid="12143" heatid="14749" lane="3" entrytime="00:01:21.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.36" />
                    <SPLIT distance="50" swimtime="00:00:37.99" />
                    <SPLIT distance="75" swimtime="00:00:58.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="426" swimtime="00:01:06.76" resultid="12144" heatid="14776" lane="4" entrytime="00:01:07.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="75" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Zürcher" birthdate="2006-12-02" gender="F" nation="SUI" license="3621" swrid="5387508" athleteid="12185">
              <RESULTS>
                <RESULT eventid="1108" points="391" swimtime="00:01:14.63" resultid="12186" heatid="14690" lane="1" entrytime="00:01:14.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.06" />
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="75" swimtime="00:00:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="347" swimtime="00:01:18.04" resultid="12187" heatid="14711" lane="4" entrytime="00:01:19.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.86" />
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="75" swimtime="00:00:58.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="487" swimtime="00:01:03.86" resultid="12188" heatid="14778" lane="4" entrytime="00:01:04.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="75" swimtime="00:00:47.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessia" lastname="Wieland" birthdate="2010-09-01" gender="F" nation="SUI" license="42277" swrid="5559295" athleteid="12176">
              <RESULTS>
                <RESULT eventid="1078" points="124" swimtime="00:01:50.01" resultid="12177" heatid="14546" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.24" />
                    <SPLIT distance="50" swimtime="00:00:51.37" />
                    <SPLIT distance="75" swimtime="00:01:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="140" swimtime="00:01:59.93" resultid="12178" heatid="14603" lane="4" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.15" />
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                    <SPLIT distance="75" swimtime="00:01:27.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="161" swimtime="00:01:32.18" resultid="12179" heatid="14649" lane="2" entrytime="00:01:38.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.36" />
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="75" swimtime="00:01:08.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Chloé" lastname="Hersberger" birthdate="2011-04-07" gender="F" nation="SUI" license="34881" swrid="4574328" athleteid="12133">
              <RESULTS>
                <RESULT eventid="1068" points="197" swimtime="00:01:33.73" resultid="12134" heatid="14521" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.65" />
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="75" swimtime="00:01:06.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="336" swimtime="00:01:29.65" resultid="12135" heatid="14609" lane="1" entrytime="00:01:34.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.63" />
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="75" swimtime="00:01:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="310" swimtime="00:01:14.18" resultid="12136" heatid="14659" lane="4" entrytime="00:01:14.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.03" />
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                    <SPLIT distance="75" swimtime="00:00:55.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathalie" lastname="Bovier" birthdate="2007-06-25" gender="F" nation="SUI" license="3887" swrid="5242993" athleteid="12121">
              <RESULTS>
                <RESULT eventid="1114" points="403" swimtime="00:01:14.27" resultid="12122" heatid="14714" lane="4" entrytime="00:01:13.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.15" />
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                    <SPLIT distance="75" swimtime="00:00:54.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="374" swimtime="00:01:26.55" resultid="12123" heatid="14747" lane="3" entrytime="00:01:26.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.94" />
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="75" swimtime="00:01:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="498" swimtime="00:01:03.37" resultid="12124" heatid="14779" lane="3" entrytime="00:01:03.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.94" />
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="75" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana Maria" lastname="Biehl" birthdate="2011-09-01" gender="F" nation="SUI" license="42276" swrid="5559907" athleteid="12113">
              <RESULTS>
                <RESULT eventid="1078" points="166" swimtime="00:01:39.69" resultid="12114" heatid="14546" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.75" />
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="75" swimtime="00:01:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="156" swimtime="00:01:55.79" resultid="12115" heatid="14603" lane="1" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.24" />
                    <SPLIT distance="50" swimtime="00:00:54.45" />
                    <SPLIT distance="75" swimtime="00:01:25.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="150" swimtime="00:01:34.50" resultid="12116" heatid="14648" lane="1" entrytime="00:01:41.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                    <SPLIT distance="75" swimtime="00:01:09.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="488" swimtime="00:02:10.01" resultid="12189" heatid="14733" lane="4" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="75" swimtime="00:00:50.19" />
                    <SPLIT distance="100" swimtime="00:01:09.88" />
                    <SPLIT distance="125" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:01:41.41" />
                    <SPLIT distance="175" swimtime="00:01:55.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12121" number="1" />
                    <RELAYPOSITION athleteid="12141" number="2" />
                    <RELAYPOSITION athleteid="12185" number="3" />
                    <RELAYPOSITION athleteid="12164" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer 3) (Zeit: 11:15)" eventid="1084" status="DSQ" swimtime="00:02:26.01" resultid="12190" heatid="14580" lane="4" entrytime="00:02:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.68" />
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="75" swimtime="00:00:57.54" />
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                    <SPLIT distance="125" swimtime="00:01:34.59" />
                    <SPLIT distance="150" swimtime="00:01:52.58" />
                    <SPLIT distance="175" swimtime="00:02:08.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12113" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="12176" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="12117" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="12133" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BREM" nation="SUI" region="RZO" clubid="12857" swrid="65617" name="SC Region Bremgarten" shortname="Brem">
          <ATHLETES>
            <ATHLETE firstname="Liun" lastname="Metzger" birthdate="2010-06-04" gender="M" nation="SUI" license="122871" swrid="5387431" athleteid="12902">
              <RESULTS>
                <RESULT eventid="1081" points="186" swimtime="00:01:24.66" resultid="12903" heatid="14558" lane="3">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.50" />
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="75" swimtime="00:01:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="212" swimtime="00:01:32.80" resultid="12904" heatid="14629" lane="4" entrytime="00:01:33.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.21" />
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                    <SPLIT distance="75" swimtime="00:01:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="236" swimtime="00:01:12.71" resultid="12905" heatid="14680" lane="2" entrytime="00:01:14.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.66" />
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="75" swimtime="00:00:55.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noah" lastname="Roth" birthdate="2007-11-03" gender="M" nation="SUI" license="114199" swrid="5227823" athleteid="12906">
              <RESULTS>
                <RESULT eventid="1117" points="254" swimtime="00:01:16.30" resultid="12907" heatid="14724" lane="4" entrytime="00:01:17.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.22" />
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="75" swimtime="00:00:56.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="313" swimtime="00:01:06.18" resultid="12908" heatid="14788" lane="2" entrytime="00:01:08.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.82" />
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="75" swimtime="00:00:49.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Wartmann" birthdate="2010-08-11" gender="F" nation="SUI" license="120487" swrid="5337119" athleteid="12919">
              <RESULTS>
                <RESULT eventid="1078" points="317" swimtime="00:01:20.45" resultid="12920" heatid="14553" lane="4" entrytime="00:01:23.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.35" />
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="75" swimtime="00:01:00.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="316" swimtime="00:01:31.46" resultid="12921" heatid="14610" lane="4" entrytime="00:01:30.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.13" />
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="75" swimtime="00:01:07.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="318" swimtime="00:01:13.58" resultid="12922" heatid="14660" lane="3" entrytime="00:01:12.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.78" />
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="75" swimtime="00:00:55.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luca" lastname="Stutz" birthdate="2007-10-11" gender="M" nation="SUI" license="2324586" swrid="4941079" athleteid="12916">
              <RESULTS>
                <RESULT eventid="1117" points="307" swimtime="00:01:11.64" resultid="12917" heatid="14726" lane="4" entrytime="00:01:11.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="75" swimtime="00:00:53.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="436" swimtime="00:00:59.23" resultid="12918" heatid="14793" lane="2" entrytime="00:00:59.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.37" />
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="75" swimtime="00:00:44.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabia" lastname="Koch" birthdate="2007-07-27" gender="F" nation="SUI" license="109775" swrid="5168000" athleteid="12878">
              <RESULTS>
                <RESULT eventid="1108" points="406" swimtime="00:01:13.71" resultid="12879" heatid="14689" lane="2" entrytime="00:01:15.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.20" />
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="75" swimtime="00:00:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="338" swimtime="00:01:18.79" resultid="12880" heatid="14711" lane="1" entrytime="00:01:18.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.24" />
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="75" swimtime="00:00:59.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="465" swimtime="00:01:04.86" resultid="12881" heatid="14778" lane="1" entrytime="00:01:04.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.88" />
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="75" swimtime="00:00:48.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amely" lastname="Manz" birthdate="2011-10-10" gender="F" nation="SUI" license="122839" swrid="5382266" athleteid="12882">
              <RESULTS>
                <RESULT eventid="1068" points="163" swimtime="00:01:39.94" resultid="12883" heatid="14520" lane="3" entrytime="00:01:40.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.52" />
                    <SPLIT distance="50" swimtime="00:00:44.31" />
                    <SPLIT distance="75" swimtime="00:01:12.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="256" swimtime="00:01:26.43" resultid="12884" heatid="14551" lane="2" entrytime="00:01:34.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.87" />
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="333" swimtime="00:01:12.46" resultid="12885" heatid="14659" lane="3" entrytime="00:01:14.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.81" />
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="75" swimtime="00:00:54.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tys" lastname="Brouwers" birthdate="2010-01-24" gender="M" nation="SUI" license="2302776" swrid="4531629" athleteid="12862">
              <RESULTS>
                <RESULT eventid="1081" points="185" swimtime="00:01:24.79" resultid="12863" heatid="14570" lane="3" entrytime="00:01:36.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.39" />
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="190" swimtime="00:01:36.15" resultid="12864" heatid="14627" lane="2" entrytime="00:01:41.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.55" />
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                    <SPLIT distance="75" swimtime="00:01:10.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 14:46)" eventid="1105" status="DSQ" swimtime="00:01:22.77" resultid="12865" heatid="14675" lane="2" entrytime="00:01:31.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.38" />
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                    <SPLIT distance="75" swimtime="00:01:01.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jamiro" lastname="Santoro" birthdate="2011-05-11" gender="M" nation="SUI" license="1772935" swrid="5466233" athleteid="12909">
              <RESULTS>
                <RESULT eventid="1081" points="86" swimtime="00:01:49.43" resultid="12910" heatid="14564" lane="1" entrytime="00:01:56.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.78" />
                    <SPLIT distance="50" swimtime="00:00:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="86" swimtime="00:01:41.52" resultid="12911" heatid="14669" lane="2" entrytime="00:01:49.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vivien" lastname="Schürch" birthdate="2011-06-10" gender="F" nation="SUI" license="124798" swrid="5426748" athleteid="12912">
              <RESULTS>
                <RESULT eventid="1078" points="183" swimtime="00:01:36.64" resultid="12913" heatid="14545" lane="4" entrytime="00:01:46.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.15" />
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="253" swimtime="00:01:38.59" resultid="12914" heatid="14605" lane="3" entrytime="00:01:45.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.76" />
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="207" swimtime="00:01:24.91" resultid="12915" heatid="14654" lane="4" entrytime="00:01:26.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.77" />
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                    <SPLIT distance="75" swimtime="00:01:03.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Fischer" birthdate="2008-01-22" gender="M" nation="GER" license="111557" swrid="4627632" athleteid="12874">
              <RESULTS>
                <RESULT eventid="1117" points="261" swimtime="00:01:15.62" resultid="12875" heatid="14723" lane="3" entrytime="00:01:19.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.96" />
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="75" swimtime="00:00:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="280" swimtime="00:01:24.58" resultid="12876" heatid="14758" lane="1" entrytime="00:01:27.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="75" swimtime="00:01:02.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="314" swimtime="00:01:06.10" resultid="12877" heatid="14788" lane="1" entrytime="00:01:09.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                    <SPLIT distance="75" swimtime="00:00:49.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mike" lastname="Wartmann" birthdate="2012-09-05" gender="M" nation="SUI" license="1772390" swrid="5440452" athleteid="12927">
              <RESULTS>
                <RESULT eventid="1081" points="156" swimtime="00:01:29.59" resultid="12928" heatid="14558" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.22" />
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="75" swimtime="00:01:06.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="144" swimtime="00:01:45.43" resultid="12929" heatid="14614" lane="1">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.39" />
                    <SPLIT distance="50" swimtime="00:00:51.07" />
                    <SPLIT distance="75" swimtime="00:01:18.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="185" swimtime="00:01:18.73" resultid="12930" heatid="14678" lane="2" entrytime="00:01:22.14">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.14" />
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="75" swimtime="00:00:59.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilia" lastname="Bellia" birthdate="2009-10-18" gender="F" nation="SUI" license="1799720" swrid="5467957" athleteid="12858">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="12859" entrytime="00:01:31.17" entrycourse="SCM" />
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="12860" entrytime="00:01:27.25" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="12861" entrytime="00:01:14.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jasper" lastname="Matter" birthdate="2010-07-27" gender="M" nation="SUI" license="1720247" swrid="5439447" athleteid="12894">
              <RESULTS>
                <RESULT eventid="1081" points="163" swimtime="00:01:28.32" resultid="12895" heatid="14571" lane="3" entrytime="00:01:31.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.22" />
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="75" swimtime="00:01:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="166" swimtime="00:01:40.62" resultid="12896" heatid="14627" lane="4" entrytime="00:01:43.84">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.70" />
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                    <SPLIT distance="75" swimtime="00:01:13.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="207" swimtime="00:01:15.94" resultid="12897" heatid="14679" lane="4" entrytime="00:01:22.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.64" />
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="75" swimtime="00:00:57.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Szonja" lastname="Merenyi" birthdate="2011-06-06" gender="F" nation="HUN" license="32635" swrid="5467960" athleteid="12898">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="12899" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="12900" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="12901" entrytime="00:01:35.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Zbinden" birthdate="2010-02-27" gender="F" nation="SUI" license="121766" swrid="5353379" athleteid="12931">
              <RESULTS>
                <RESULT eventid="1078" points="214" swimtime="00:01:31.64" resultid="12932" heatid="14552" lane="1" entrytime="00:01:33.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.74" />
                    <SPLIT distance="50" swimtime="00:00:44.70" />
                    <SPLIT distance="75" swimtime="00:01:09.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="285" swimtime="00:01:34.73" resultid="12933" heatid="14609" lane="4" entrytime="00:01:34.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                    <SPLIT distance="75" swimtime="00:01:10.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="279" swimtime="00:01:16.86" resultid="12934" heatid="14658" lane="3" entrytime="00:01:20.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.18" />
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="75" swimtime="00:00:57.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liv" lastname="Martin" birthdate="2010-01-09" gender="F" nation="SUI" license="1772928" swrid="5442079" athleteid="12890">
              <RESULTS>
                <RESULT eventid="1078" status="DNS" swimtime="00:00:00.00" resultid="12891" heatid="14552" lane="2" entrytime="00:01:24.00" />
                <RESULT eventid="1092" points="420" swimtime="00:01:23.27" resultid="12892" heatid="14610" lane="2" entrytime="00:01:23.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                    <SPLIT distance="75" swimtime="00:01:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="448" swimtime="00:01:05.64" resultid="12893" heatid="14661" lane="3" entrytime="00:01:08.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="75" swimtime="00:00:48.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ronja" lastname="Dobler" birthdate="2006-10-07" gender="F" nation="SUI" license="109777" swrid="5167985" athleteid="12870">
              <RESULTS>
                <RESULT eventid="1108" points="403" swimtime="00:01:13.93" resultid="12871" heatid="14691" lane="3" entrytime="00:01:11.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.03" />
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="75" swimtime="00:00:54.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="414" swimtime="00:01:13.59" resultid="12872" heatid="14713" lane="3" entrytime="00:01:14.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.24" />
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="75" swimtime="00:00:54.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="411" swimtime="00:01:07.58" resultid="12873" heatid="14777" lane="1" entrytime="00:01:05.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.29" />
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="75" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessio" lastname="Chechele" birthdate="2008-08-21" gender="M" nation="SUI" license="2310645" swrid="4941100" athleteid="12866">
              <RESULTS>
                <RESULT eventid="1117" points="218" swimtime="00:01:20.23" resultid="12867" heatid="14722" lane="1" entrytime="00:01:24.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.44" />
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="75" swimtime="00:01:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="233" swimtime="00:01:29.87" resultid="12868" heatid="14757" lane="3" entrytime="00:01:29.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.64" />
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="75" swimtime="00:01:06.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="308" swimtime="00:01:06.54" resultid="12869" heatid="14788" lane="3" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.98" />
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="75" swimtime="00:00:49.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ava" lastname="Martin" birthdate="2008-03-03" gender="F" nation="SUI" license="1772925" swrid="5442078" athleteid="12886">
              <RESULTS>
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="12887" entrytime="00:01:27.21" entrycourse="SCM" />
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="12888" entrytime="00:01:28.32" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="12889" entrytime="00:01:14.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucy" lastname="Wartmann" birthdate="2007-01-11" gender="F" nation="SUI" license="110236" swrid="5185893" athleteid="12923">
              <RESULTS>
                <RESULT eventid="1114" points="377" swimtime="00:01:15.95" resultid="12924" heatid="14713" lane="1" entrytime="00:01:15.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.98" />
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="75" swimtime="00:00:56.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="317" swimtime="00:01:31.45" resultid="12925" heatid="14744" lane="1" entrytime="00:01:31.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.35" />
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                    <SPLIT distance="75" swimtime="00:01:07.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="335" swimtime="00:01:12.34" resultid="12926" heatid="14773" lane="3" entrytime="00:01:10.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="75" swimtime="00:00:53.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="194" swimtime="00:02:21.07" resultid="12935" heatid="14818" lane="4" entrytime="00:02:25.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:53.67" />
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="75" swimtime="00:01:29.58" />
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                    <SPLIT distance="125" swimtime="00:02:04.16" />
                    <SPLIT distance="150" swimtime="00:01:48.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12894" number="1" />
                    <RELAYPOSITION athleteid="12927" number="2" />
                    <RELAYPOSITION athleteid="12862" number="3" />
                    <RELAYPOSITION athleteid="12902" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="290" swimtime="00:02:16.63" resultid="12936" heatid="14735" lane="3" entrytime="00:02:25.77">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.68" />
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="75" swimtime="00:00:52.92" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="125" swimtime="00:01:31.14" />
                    <SPLIT distance="150" swimtime="00:01:50.59" />
                    <SPLIT distance="175" swimtime="00:02:03.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12866" number="1" />
                    <RELAYPOSITION athleteid="12906" number="2" />
                    <RELAYPOSITION athleteid="12874" number="3" />
                    <RELAYPOSITION athleteid="12916" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="292" swimtime="00:02:19.29" resultid="12937" heatid="14817" lane="1" entrytime="00:02:18.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.21" />
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="75" swimtime="00:00:53.46" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="125" swimtime="00:01:28.44" />
                    <SPLIT distance="150" swimtime="00:01:45.52" />
                    <SPLIT distance="175" swimtime="00:02:01.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12931" number="1" />
                    <RELAYPOSITION athleteid="12912" number="2" />
                    <RELAYPOSITION athleteid="12919" number="3" />
                    <RELAYPOSITION athleteid="12882" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" status="WDR" swimtime="00:00:00.00" resultid="12938" entrytime="00:02:17.84">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12923" number="1" />
                    <RELAYPOSITION athleteid="12858" number="2" />
                    <RELAYPOSITION athleteid="12878" number="3" />
                    <RELAYPOSITION athleteid="12870" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="AARE" nation="SUI" region="RZW" clubid="12199" swrid="65609" name="Schwimmclub Aarefisch Aarau" shortname="Schwimmclub Aarefisch">
          <ATHLETES>
            <ATHLETE firstname="Miro" lastname="Hunziker" birthdate="2012-11-22" gender="M" nation="SUI" license="31957" swrid="5464171" athleteid="14093">
              <RESULTS>
                <RESULT eventid="1081" points="100" swimtime="00:01:43.90" resultid="14094" heatid="14565" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.59" />
                    <SPLIT distance="50" swimtime="00:00:49.45" />
                    <SPLIT distance="75" swimtime="00:01:17.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="91" swimtime="00:02:02.63" resultid="14095" heatid="14621" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.51" />
                    <SPLIT distance="75" swimtime="00:01:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="96" swimtime="00:01:37.83" resultid="14096" heatid="14670" lane="1" entrytime="00:01:47.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.87" />
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="75" swimtime="00:01:12.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michelle" lastname="Saxer" birthdate="2007-02-17" gender="F" nation="SUI" license="24849" swrid="4995456" athleteid="14217">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="14218" entrytime="00:01:15.77" entrycourse="SCM" />
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="14219" entrytime="00:01:16.85" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="14220" entrytime="00:01:09.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maxime" lastname="Kiliçer" birthdate="2011-07-06" gender="M" nation="SUI" swrid="5551356" athleteid="14112">
              <RESULTS>
                <RESULT eventid="1081" points="74" swimtime="00:01:54.67" resultid="14113" heatid="14560" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.95" />
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                    <SPLIT distance="75" swimtime="00:01:25.15" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...) (Zeit: 12:45)" eventid="1095" status="DSQ" swimtime="00:02:12.76" resultid="14114" heatid="14615" lane="3" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.32" />
                    <SPLIT distance="50" swimtime="00:01:02.77" />
                    <SPLIT distance="75" swimtime="00:01:37.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="97" swimtime="00:01:37.55" resultid="14115" heatid="14667" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.03" />
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jonathan" lastname="Thölking" birthdate="2015-01-09" gender="M" nation="SUI" athleteid="14257">
              <RESULTS>
                <RESULT eventid="1076" points="51" swimtime="00:00:59.74" resultid="14258" heatid="14534" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="527 - Wechselbeinschlag während des Schwimmens (Zeit: 11:54)" eventid="1090" status="DSQ" swimtime="00:01:25.22" resultid="14259" heatid="14591" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 13:30)" eventid="1100" status="DSQ" swimtime="00:00:58.29" resultid="14260" heatid="14638" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yannick" lastname="Rohr" birthdate="2006-12-05" gender="M" nation="SUI" license="24916" swrid="5257642" athleteid="14202">
              <RESULTS>
                <RESULT eventid="1111" points="313" swimtime="00:01:10.32" resultid="14203" heatid="14697" lane="2" entrytime="00:01:12.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.99" />
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="75" swimtime="00:00:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="289" swimtime="00:01:13.04" resultid="14204" heatid="14725" lane="3" entrytime="00:01:12.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.57" />
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="75" swimtime="00:00:53.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="296" swimtime="00:01:22.97" resultid="14205" heatid="14759" lane="1" entrytime="00:01:24.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.41" />
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                    <SPLIT distance="75" swimtime="00:01:01.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="377" swimtime="00:01:02.17" resultid="14206" heatid="14792" lane="4" entrytime="00:01:01.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.60" />
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="75" swimtime="00:00:45.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danyal" lastname="Nisamov" birthdate="2010-07-18" gender="M" nation="SUI" license="24754" swrid="5329310" athleteid="14163">
              <RESULTS>
                <RESULT eventid="1071" points="81" swimtime="00:01:50.33" resultid="14164" heatid="14523" lane="1" entrytime="00:02:21.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.36" />
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                    <SPLIT distance="75" swimtime="00:01:19.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="179" swimtime="00:01:25.75" resultid="14165" heatid="14572" lane="2" entrytime="00:01:28.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.17" />
                    <SPLIT distance="50" swimtime="00:00:41.76" />
                    <SPLIT distance="75" swimtime="00:01:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="165" swimtime="00:01:40.78" resultid="14166" heatid="14626" lane="1" entrytime="00:01:47.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.99" />
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                    <SPLIT distance="75" swimtime="00:01:14.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 14:55)" eventid="1105" status="DSQ" swimtime="00:01:14.94" resultid="14167" heatid="14680" lane="4" entrytime="00:01:17.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="75" swimtime="00:00:55.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Thölking" birthdate="2009-09-04" gender="M" nation="SUI" license="24807" swrid="5159306" athleteid="14261">
              <RESULTS>
                <RESULT eventid="1111" points="302" swimtime="00:01:11.17" resultid="14262" heatid="14697" lane="3" entrytime="00:01:15.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.22" />
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="75" swimtime="00:00:51.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="312" swimtime="00:01:11.24" resultid="14263" heatid="14727" lane="1" entrytime="00:01:09.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.17" />
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="75" swimtime="00:00:53.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="298" swimtime="00:01:22.76" resultid="14264" heatid="14759" lane="4" entrytime="00:01:25.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                    <SPLIT distance="75" swimtime="00:01:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="404" swimtime="00:01:00.78" resultid="14265" heatid="14793" lane="3" entrytime="00:00:59.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.61" />
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="75" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hordi" lastname="Konaschenkov" birthdate="2012-02-29" gender="M" nation="UKR" license="42614" athleteid="14116">
              <RESULTS>
                <RESULT eventid="1081" points="102" swimtime="00:01:43.36" resultid="14117" heatid="14563" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.09" />
                    <SPLIT distance="75" swimtime="00:01:18.14" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  2) (Zeit: 12:54)" eventid="1095" status="DSQ" swimtime="00:01:56.22" resultid="14118" heatid="14618" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.88" />
                    <SPLIT distance="50" swimtime="00:00:54.21" />
                    <SPLIT distance="75" swimtime="00:01:26.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="129" swimtime="00:01:28.92" resultid="14119" heatid="14669" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.95" />
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                    <SPLIT distance="75" swimtime="00:01:08.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lars" lastname="Oeschger" birthdate="2007-09-11" gender="M" nation="SUI" license="24819" swrid="5159319" athleteid="14173">
              <RESULTS>
                <RESULT eventid="1111" points="357" swimtime="00:01:07.31" resultid="14174" heatid="14699" lane="4" entrytime="00:01:07.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.23" />
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                    <SPLIT distance="75" swimtime="00:00:48.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="268" swimtime="00:01:14.88" resultid="14175" heatid="14724" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.97" />
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                    <SPLIT distance="75" swimtime="00:00:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="294" swimtime="00:01:23.22" resultid="14176" heatid="14757" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.83" />
                    <SPLIT distance="50" swimtime="00:00:38.55" />
                    <SPLIT distance="75" swimtime="00:01:00.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="394" swimtime="00:01:01.26" resultid="14177" heatid="14791" lane="3" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.12" />
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="75" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luc Joël" lastname="Nef" birthdate="2010-09-15" gender="M" nation="SUI" license="25086" swrid="5440234" athleteid="14152">
              <RESULTS>
                <RESULT eventid="1081" points="64" swimtime="00:02:00.37" resultid="14153" heatid="14561" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.41" />
                    <SPLIT distance="50" swimtime="00:00:55.10" />
                    <SPLIT distance="75" swimtime="00:01:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="37" swimtime="00:02:45.55" resultid="14154" heatid="14617" lane="4" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.71" />
                    <SPLIT distance="50" swimtime="00:01:15.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="65" swimtime="00:01:51.46" resultid="14155" heatid="14667" lane="1" entrytime="00:02:01.82">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.30" />
                    <SPLIT distance="50" swimtime="00:00:50.21" />
                    <SPLIT distance="75" swimtime="00:01:20.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Twyla" lastname="Reinhard" birthdate="2005-10-09" gender="F" nation="SUI" license="19736" swrid="5104838" athleteid="14192">
              <RESULTS>
                <RESULT eventid="1108" points="543" swimtime="00:01:06.90" resultid="14193" heatid="14692" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="75" swimtime="00:00:48.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="552" swimtime="00:01:06.91" resultid="14194" heatid="14716" lane="4" entrytime="00:01:06.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="75" swimtime="00:00:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="431" swimtime="00:01:22.55" resultid="14195" heatid="14748" lane="1" entrytime="00:01:24.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.57" />
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="75" swimtime="00:01:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="583" swimtime="00:01:00.15" resultid="14196" heatid="14781" lane="1" entrytime="00:00:59.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.74" />
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                    <SPLIT distance="75" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="579" swimtime="00:00:30.71" resultid="14846" heatid="14801" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6681" points="452" swimtime="00:00:37.21" resultid="14863" heatid="14803" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6635" points="501" swimtime="00:00:30.69" resultid="14872" heatid="14805" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilie" lastname="Sandberg" birthdate="2011-05-16" gender="F" nation="SWE" license="24768" swrid="5043646" athleteid="14212">
              <RESULTS>
                <RESULT eventid="1068" points="96" swimtime="00:01:59.04" resultid="14213" heatid="14517" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:26.44" />
                    <SPLIT distance="50" swimtime="00:00:54.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="189" swimtime="00:01:35.64" resultid="14214" heatid="14550" lane="4" entrytime="00:01:36.53">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.30" />
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="75" swimtime="00:01:11.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="171" swimtime="00:01:52.22" resultid="14215" heatid="14600" lane="3" entrytime="00:02:02.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.67" />
                    <SPLIT distance="50" swimtime="00:00:53.39" />
                    <SPLIT distance="75" swimtime="00:01:22.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="241" swimtime="00:01:20.71" resultid="14216" heatid="14657" lane="3" entrytime="00:01:22.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.00" />
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="75" swimtime="00:01:00.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Chiara" lastname="Haller" birthdate="2007-01-01" gender="F" nation="SUI" swrid="4889154" athleteid="14076">
              <RESULTS>
                <RESULT eventid="1108" points="483" swimtime="00:01:09.56" resultid="14077" heatid="14691" lane="1" entrytime="00:01:12.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="75" swimtime="00:00:50.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="437" swimtime="00:01:12.28" resultid="14078" heatid="14715" lane="4" entrytime="00:01:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.47" />
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="75" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="557" swimtime="00:01:15.77" resultid="14079" heatid="14749" lane="2" entrytime="00:01:16.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.31" />
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="75" swimtime="00:00:55.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="546" swimtime="00:01:01.45" resultid="14080" heatid="14779" lane="1" entrytime="00:01:03.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.24" />
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="75" swimtime="00:00:45.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="431" swimtime="00:00:33.88" resultid="14848" heatid="14842" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sven" lastname="Thalmann" birthdate="1999-08-21" gender="M" nation="SUI" license="24904" swrid="4233857" athleteid="14252">
              <RESULTS>
                <RESULT eventid="1111" points="383" swimtime="00:01:05.76" resultid="14253" heatid="14700" lane="3" entrytime="00:01:03.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="75" swimtime="00:00:48.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="390" swimtime="00:01:06.11" resultid="14254" heatid="14729" lane="4" entrytime="00:01:04.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="75" swimtime="00:00:49.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="376" swimtime="00:01:16.65" resultid="14255" heatid="14762" lane="1" entrytime="00:01:12.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.74" />
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="75" swimtime="00:00:56.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="464" swimtime="00:00:58.03" resultid="14256" heatid="14795" lane="4" entrytime="00:00:57.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.68" />
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nadine" lastname="Haas" birthdate="2009-10-27" gender="F" nation="SUI" swrid="5503632" athleteid="14072">
              <RESULTS>
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="14073" entrytime="00:01:45.00" />
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="14074" entrytime="00:02:00.00" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="14075" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malte" lastname="Rohden" birthdate="1995-09-28" gender="M" nation="GER" license="25142" swrid="4666668" athleteid="14197">
              <RESULTS>
                <RESULT eventid="1111" points="430" swimtime="00:01:03.30" resultid="14198" heatid="14700" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="75" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="450" swimtime="00:01:03.05" resultid="14199" heatid="14729" lane="1" entrytime="00:01:04.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="75" swimtime="00:00:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="497" swimtime="00:01:09.86" resultid="14200" heatid="14763" lane="1" entrytime="00:01:05.71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="75" swimtime="00:00:51.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="508" swimtime="00:00:56.29" resultid="14201" heatid="14794" lane="2" entrytime="00:00:58.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.89" />
                    <SPLIT distance="50" swimtime="00:00:26.92" />
                    <SPLIT distance="75" swimtime="00:00:41.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Morini" birthdate="2006-07-10" gender="F" nation="SUI" license="24786" swrid="5103076" athleteid="14139">
              <RESULTS>
                <RESULT eventid="1108" points="271" swimtime="00:01:24.37" resultid="14140" heatid="14689" lane="4" entrytime="00:01:20.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.16" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:01:00.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="367" swimtime="00:01:16.61" resultid="14141" heatid="14712" lane="3" entrytime="00:01:17.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.40" />
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="75" swimtime="00:00:57.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="361" swimtime="00:01:10.55" resultid="14142" heatid="14776" lane="3" entrytime="00:01:06.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="75" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natascha" lastname="Stucki" birthdate="2013-05-10" gender="F" nation="SUI" license="29573" swrid="5456696" athleteid="14234">
              <RESULTS>
                <RESULT eventid="1064" points="73" swimtime="00:00:58.19" resultid="14235" heatid="14513" lane="3" entrytime="00:01:00.49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="103" swimtime="00:00:54.50" resultid="14236" heatid="14532" lane="1" entrytime="00:00:54.75">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="84" swimtime="00:01:05.10" resultid="14237" heatid="14585" lane="3" entrytime="00:01:17.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="119" swimtime="00:00:46.49" resultid="14238" heatid="14636" lane="4" entrytime="00:00:48.79">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kian" lastname="Pourtehrani" birthdate="2011-07-03" gender="M" nation="SUI" license="25092" swrid="5382270" athleteid="14178">
              <RESULTS>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 10:25)" eventid="1081" status="DSQ" swimtime="00:01:40.70" resultid="14179" heatid="14562" lane="2" entrytime="00:02:01.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.94" />
                    <SPLIT distance="50" swimtime="00:00:51.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="90" swimtime="00:02:03.37" resultid="14180" heatid="14616" lane="2" entrytime="00:02:23.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.66" />
                    <SPLIT distance="50" swimtime="00:00:57.62" />
                    <SPLIT distance="75" swimtime="00:01:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="139" swimtime="00:01:26.65" resultid="14181" heatid="14674" lane="1" entrytime="00:01:33.91">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="75" swimtime="00:01:05.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline Zoé" lastname="Nef" birthdate="2014-07-14" gender="F" nation="SUI" swrid="5538024" athleteid="14148">
              <RESULTS>
                <RESULT eventid="1074" points="42" swimtime="00:01:13.62" resultid="14149" heatid="14527" lane="1" entrytime="00:01:20.42">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="33" swimtime="00:01:28.69" resultid="14150" heatid="14584" lane="4" entrytime="00:01:45.27" />
                <RESULT eventid="1098" points="22" swimtime="00:01:21.59" resultid="14151" heatid="14631" lane="1" entrytime="00:01:20.63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mailin" lastname="Hösli" birthdate="2007-07-24" gender="F" nation="SUI" license="24832" swrid="5257619" athleteid="14090">
              <RESULTS>
                <RESULT eventid="1114" points="262" swimtime="00:01:25.69" resultid="14091" heatid="14708" lane="4" entrytime="00:01:25.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.61" />
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="75" swimtime="00:01:03.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="288" swimtime="00:01:34.42" resultid="14092" heatid="14742" lane="1" entrytime="00:01:35.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                    <SPLIT distance="50" swimtime="00:00:44.58" />
                    <SPLIT distance="75" swimtime="00:01:09.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksim" lastname="Bucher" birthdate="2013-04-16" gender="M" nation="SUI" license="25085" swrid="5411014" athleteid="14027">
              <RESULTS>
                <RESULT eventid="1066" points="90" swimtime="00:00:48.48" resultid="14028" heatid="14516" lane="3" entrytime="00:01:01.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="123" swimtime="00:00:44.56" resultid="14029" heatid="14537" lane="1" entrytime="00:00:52.49">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="115" swimtime="00:00:51.85" resultid="14030" heatid="14594" lane="3" entrytime="00:00:54.98">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="160" swimtime="00:00:37.06" resultid="14031" heatid="14641" lane="2" entrytime="00:00:38.66">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samira" lastname="Arnold" birthdate="2002-04-11" gender="F" nation="SUI" license="24887" swrid="4705701" athleteid="14008">
              <RESULTS>
                <RESULT eventid="1124" points="550" swimtime="00:01:16.10" resultid="14009" heatid="14750" lane="1" entrytime="00:01:14.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.41" />
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                    <SPLIT distance="75" swimtime="00:00:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="501" swimtime="00:01:03.26" resultid="14288" heatid="14779" lane="2" entrytime="00:01:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.11" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:47.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="431" swimtime="00:00:33.87" resultid="14851" heatid="14842" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Balliello" birthdate="2008-10-28" gender="F" nation="GER" license="25082" swrid="5382274" athleteid="14011">
              <RESULTS>
                <RESULT eventid="1114" points="250" swimtime="00:01:27.08" resultid="14012" heatid="14706" lane="1" entrytime="00:01:30.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="75" swimtime="00:01:05.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="284" swimtime="00:01:34.86" resultid="14013" heatid="14741" lane="2" entrytime="00:01:37.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.96" />
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="75" swimtime="00:01:10.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriele" lastname="Marinucci" birthdate="2004-01-03" gender="M" nation="SUI" license="24783" swrid="4964846" athleteid="14129">
              <RESULTS>
                <RESULT eventid="1117" status="WDR" swimtime="00:00:00.00" resultid="14130" entrytime="00:01:00.91" entrycourse="SCM" />
                <RESULT eventid="1127" status="WDR" swimtime="00:00:00.00" resultid="14131" entrytime="00:01:11.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noemi" lastname="Maurer" birthdate="2013-04-02" gender="F" nation="SUI" swrid="5481978" athleteid="14132">
              <RESULTS>
                <RESULT eventid="1074" points="93" swimtime="00:00:56.42" resultid="14133" heatid="14529" lane="2" entrytime="00:01:02.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="75" swimtime="00:01:07.71" resultid="14134" heatid="14586" lane="1" entrytime="00:01:11.56">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="80" swimtime="00:00:53.20" resultid="14135" heatid="14634" lane="1" entrytime="00:00:57.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fiona" lastname="Weber" birthdate="2013-07-25" gender="F" nation="SUI" swrid="5489045" athleteid="14271">
              <RESULTS>
                <RESULT eventid="1074" points="58" swimtime="00:01:06.10" resultid="14272" heatid="14528" lane="1" entrytime="00:01:11.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="55" swimtime="00:01:14.84" resultid="14273" heatid="14585" lane="4" entrytime="00:01:19.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="46" swimtime="00:01:03.84" resultid="14274" heatid="14631" lane="3" entrytime="00:01:14.64" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jens" lastname="Oeschger" birthdate="2010-09-19" gender="M" nation="SUI" license="24803" swrid="5302397" athleteid="14168">
              <RESULTS>
                <RESULT eventid="1071" points="195" swimtime="00:01:22.35" resultid="14169" heatid="14526" lane="4" entrytime="00:01:26.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="75" swimtime="00:00:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="203" swimtime="00:01:22.21" resultid="14170" heatid="14573" lane="4" entrytime="00:01:24.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.10" />
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                    <SPLIT distance="75" swimtime="00:01:01.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="141" swimtime="00:01:46.20" resultid="14171" heatid="14623" lane="2" entrytime="00:01:52.81">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.88" />
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="75" swimtime="00:01:17.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="249" swimtime="00:01:11.39" resultid="14172" heatid="14681" lane="1" entrytime="00:01:12.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.39" />
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="75" swimtime="00:00:53.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Hauss" birthdate="2014-10-10" gender="M" nation="SUI" license="34379" swrid="5509057" athleteid="14081">
              <RESULTS>
                <RESULT eventid="1076" points="69" swimtime="00:00:54.05" resultid="14082" heatid="14536" lane="3" entrytime="00:00:58.38">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="69" swimtime="00:01:01.43" resultid="14083" heatid="14593" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="86" swimtime="00:00:45.53" resultid="14084" heatid="14640" lane="3" entrytime="00:00:49.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Añón" birthdate="2013-05-21" gender="F" nation="SUI" license="29352" swrid="5456690" athleteid="13998">
              <RESULTS>
                <RESULT eventid="1064" points="52" swimtime="00:01:05.00" resultid="13999" heatid="14513" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="84" swimtime="00:00:58.23" resultid="14000" heatid="14531" lane="2" entrytime="00:00:58.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="93" swimtime="00:01:02.82" resultid="14001" heatid="14586" lane="3" entrytime="00:01:10.61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="61" swimtime="00:00:58.07" resultid="14002" heatid="14633" lane="3" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Hofmann" birthdate="2007-02-14" gender="M" nation="SUI" license="24717" swrid="4889163" athleteid="14085">
              <RESULTS>
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="14086" entrytime="00:01:17.31" entrycourse="SCM" />
                <RESULT eventid="1117" status="WDR" swimtime="00:00:00.00" resultid="14087" entrytime="00:01:25.00" />
                <RESULT eventid="1127" status="WDR" swimtime="00:00:00.00" resultid="14088" entrytime="00:01:25.42" entrycourse="SCM" />
                <RESULT eventid="1133" status="WDR" swimtime="00:00:00.00" resultid="14089" entrytime="00:01:01.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nino" lastname="Tahedl" birthdate="2011-09-12" gender="M" nation="SUI" license="25107" swrid="5440236" athleteid="14248">
              <RESULTS>
                <RESULT eventid="1081" points="45" swimtime="00:02:15.83" resultid="14249" heatid="14562" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.92" />
                    <SPLIT distance="50" swimtime="00:01:02.92" />
                    <SPLIT distance="75" swimtime="00:01:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Zeit: 12:44)" eventid="1095" status="DSQ" swimtime="00:02:18.97" resultid="14250" heatid="14615" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.09" />
                    <SPLIT distance="50" swimtime="00:01:04.48" />
                    <SPLIT distance="75" swimtime="00:01:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="36" swimtime="00:02:15.28" resultid="14251" heatid="14665" lane="3" entrytime="00:02:19.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.66" />
                    <SPLIT distance="75" swimtime="00:01:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Federico" lastname="Salghetti-Drioli" birthdate="2000-10-04" gender="M" nation="SUI" license="24779" swrid="4598611" athleteid="14207">
              <RESULTS>
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="14208" entrytime="00:01:01.17" entrycourse="SCM" />
                <RESULT eventid="1117" status="WDR" swimtime="00:00:00.00" resultid="14209" entrytime="00:01:04.14" entrycourse="SCM" />
                <RESULT eventid="1127" status="WDR" swimtime="00:00:00.00" resultid="14210" entrytime="00:01:12.25" entrycourse="SCM" />
                <RESULT eventid="1133" status="WDR" swimtime="00:00:00.00" resultid="14211" entrytime="00:00:54.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kevin" lastname="Affentranger" birthdate="2001-08-17" gender="M" nation="SUI" license="24816" swrid="4703382" athleteid="13988">
              <RESULTS>
                <RESULT eventid="1111" points="475" swimtime="00:01:01.20" resultid="13989" heatid="14701" lane="3" entrytime="00:00:57.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.86" />
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="75" swimtime="00:00:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="341" swimtime="00:01:09.15" resultid="13990" heatid="14728" lane="2" entrytime="00:01:04.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.15" />
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="75" swimtime="00:00:51.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="440" swimtime="00:01:12.74" resultid="13991" heatid="14763" lane="3" entrytime="00:01:04.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="75" swimtime="00:00:52.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="495" swimtime="00:00:56.80" resultid="13992" heatid="14797" lane="3" entrytime="00:00:52.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.96" />
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="75" swimtime="00:00:41.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noemi" lastname="Nguyen" birthdate="2008-12-31" gender="F" nation="SUI" license="24861" swrid="5382267" athleteid="14160">
              <RESULTS>
                <RESULT eventid="1124" status="SICK" swimtime="00:00:00.00" resultid="14161" entrytime="00:01:35.63" />
                <RESULT eventid="1108" status="SICK" swimtime="00:00:00.00" resultid="14162" entrytime="00:01:30.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alvaro" lastname="Garrido" birthdate="2010-10-28" gender="M" nation="SUI" swrid="5551355" athleteid="14064">
              <RESULTS>
                <RESULT eventid="1081" points="118" swimtime="00:01:38.45" resultid="14065" heatid="14569" lane="4" entrytime="00:01:41.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="128" swimtime="00:01:49.70" resultid="14066" heatid="14622" lane="4" entrytime="00:01:56.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.88" />
                    <SPLIT distance="50" swimtime="00:00:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="132" swimtime="00:01:28.13" resultid="14067" heatid="14677" lane="1" entrytime="00:01:27.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.31" />
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Colin" lastname="Glässel" birthdate="2013-03-11" gender="M" nation="SUI" swrid="5538022" athleteid="14068">
              <RESULTS>
                <RESULT eventid="1076" points="66" swimtime="00:00:54.84" resultid="14069" heatid="14535" lane="1" entrytime="00:01:04.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="72" swimtime="00:01:00.44" resultid="14070" heatid="14591" lane="2" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="39" swimtime="00:00:59.44" resultid="14071" heatid="14638" lane="2" entrytime="00:01:05.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefan Oliver" lastname="Mos" birthdate="2009-06-08" gender="M" nation="SUI" swrid="5503633" athleteid="14143">
              <RESULTS>
                <RESULT eventid="1111" points="152" swimtime="00:01:29.50" resultid="14144" heatid="14695" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.20" />
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="75" swimtime="00:01:02.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="194" swimtime="00:01:23.48" resultid="14145" heatid="14722" lane="3" entrytime="00:01:23.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                    <SPLIT distance="75" swimtime="00:01:02.46" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  1) (Zeit: 18:47)" eventid="1127" status="DSQ" swimtime="00:01:50.17" resultid="14146" heatid="14754" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.27" />
                    <SPLIT distance="50" swimtime="00:00:52.56" />
                    <SPLIT distance="75" swimtime="00:01:21.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="246" swimtime="00:01:11.68" resultid="14147" heatid="14787" lane="3" entrytime="00:01:10.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="75" swimtime="00:00:53.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nora" lastname="Wick" birthdate="2002-08-24" gender="F" nation="SUI" license="24863" swrid="4971878" athleteid="14275">
              <RESULTS>
                <RESULT eventid="1108" points="637" swimtime="00:01:03.44" resultid="14276" heatid="14692" lane="3" entrytime="00:01:02.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.04" />
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                    <SPLIT distance="75" swimtime="00:00:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="513" swimtime="00:01:08.56" resultid="14277" heatid="14716" lane="3" entrytime="00:01:05.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.85" />
                    <SPLIT distance="50" swimtime="00:00:32.43" />
                    <SPLIT distance="75" swimtime="00:00:50.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="470" swimtime="00:01:20.20" resultid="14278" heatid="14750" lane="4" entrytime="00:01:14.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="75" swimtime="00:00:58.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="615" swimtime="00:00:59.07" resultid="14279" heatid="14781" lane="2" entrytime="00:00:58.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.40" />
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                    <SPLIT distance="75" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="539" swimtime="00:00:31.45" resultid="14849" heatid="14842" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6681" points="505" swimtime="00:00:35.86" resultid="14864" heatid="14803" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6635" points="588" swimtime="00:00:29.10" resultid="14871" heatid="14805" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6637" points="637" swimtime="00:00:26.64" resultid="14877" heatid="14807" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonie" lastname="Sigg" birthdate="2014-02-22" gender="F" nation="SUI" swrid="5551358" athleteid="14225">
              <RESULTS>
                <RESULT eventid="1074" points="78" swimtime="00:00:59.75" resultid="14226" heatid="14527" lane="2" entrytime="00:01:12.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="62" swimtime="00:01:11.86" resultid="14227" heatid="14584" lane="1" entrytime="00:01:40.00" />
                <RESULT eventid="1098" points="58" swimtime="00:00:59.00" resultid="14228" heatid="14632" lane="1" entrytime="00:01:10.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Charlotte" lastname="Bieri" birthdate="2014-09-06" gender="F" nation="SUI" swrid="5551354" athleteid="14014">
              <RESULTS>
                <RESULT eventid="1074" points="73" swimtime="00:01:00.98" resultid="14015" heatid="14529" lane="3" entrytime="00:01:03.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="97" swimtime="00:01:01.98" resultid="14016" heatid="14589" lane="4" entrytime="00:00:58.48">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="74" swimtime="00:00:54.48" resultid="14017" heatid="14635" lane="1" entrytime="00:00:54.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessia" lastname="Sprecher" birthdate="2009-08-22" gender="F" nation="SUI" license="24715" swrid="5451774" athleteid="14229">
              <RESULTS>
                <RESULT eventid="1108" points="296" swimtime="00:01:21.90" resultid="14230" heatid="14688" lane="2" entrytime="00:01:21.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.43" />
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="75" swimtime="00:00:59.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="280" swimtime="00:01:23.89" resultid="14231" heatid="14709" lane="4" entrytime="00:01:22.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="75" swimtime="00:01:02.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="14232" entrytime="00:01:41.64" entrycourse="SCM" />
                <RESULT eventid="1130" points="383" swimtime="00:01:09.19" resultid="14233" heatid="14772" lane="4" entrytime="00:01:11.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.57" />
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="75" swimtime="00:00:51.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tobias" lastname="Dietiker" birthdate="2011-09-13" gender="M" nation="SUI" license="25084" swrid="5411019" athleteid="14050">
              <RESULTS>
                <RESULT eventid="1071" points="125" swimtime="00:01:35.45" resultid="14051" heatid="14524" lane="3" entrytime="00:02:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.55" />
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="75" swimtime="00:01:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="140" swimtime="00:01:32.88" resultid="14052" heatid="14570" lane="2" entrytime="00:01:33.69">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="156" swimtime="00:01:42.75" resultid="14053" heatid="14628" lane="1" entrytime="00:01:40.44">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.21" />
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="75" swimtime="00:01:16.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="173" swimtime="00:01:20.58" resultid="14054" heatid="14678" lane="3" entrytime="00:01:23.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.63" />
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luongo" birthdate="2013-05-29" gender="F" nation="SUI" license="28180" swrid="5445056" athleteid="14120">
              <RESULTS>
                <RESULT eventid="1064" points="89" swimtime="00:00:54.41" resultid="14121" heatid="14515" lane="1" entrytime="00:00:49.91">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="178" swimtime="00:00:45.45" resultid="14122" heatid="14533" lane="1" entrytime="00:00:46.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="139" swimtime="00:00:55.01" resultid="14123" heatid="14589" lane="3" entrytime="00:00:53.41">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="208" swimtime="00:00:38.64" resultid="14124" heatid="14637" lane="1" entrytime="00:00:40.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gion" lastname="Maissen" birthdate="2014-01-05" gender="M" nation="SUI" license="33711" swrid="5481976" athleteid="14125">
              <RESULTS>
                <RESULT eventid="1076" points="56" swimtime="00:00:58.04" resultid="14126" heatid="14534" lane="2" entrytime="00:01:05.28" />
                <RESULT eventid="1090" points="58" swimtime="00:01:05.08" resultid="14127" heatid="14592" lane="3" entrytime="00:01:10.74">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="58" swimtime="00:00:51.88" resultid="14128" heatid="14638" lane="3" entrytime="00:01:06.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michelle" lastname="Armandi" birthdate="2006-11-20" gender="F" nation="SUI" license="25152" swrid="5053783" athleteid="14003">
              <RESULTS>
                <RESULT eventid="1108" points="499" swimtime="00:01:08.84" resultid="14004" heatid="14692" lane="1" entrytime="00:01:07.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.38" />
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="75" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="459" swimtime="00:01:11.12" resultid="14005" heatid="14714" lane="2" entrytime="00:01:12.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.59" />
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="75" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="440" swimtime="00:01:21.93" resultid="14006" heatid="14748" lane="2" entrytime="00:01:22.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.53" />
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="75" swimtime="00:00:59.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="610" swimtime="00:00:59.22" resultid="14007" heatid="14781" lane="4" entrytime="00:00:59.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.31" />
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                    <SPLIT distance="75" swimtime="00:00:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="506" swimtime="00:00:32.12" resultid="14850" heatid="14842" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6681" points="430" swimtime="00:00:37.82" resultid="14865" heatid="14803" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jann" lastname="Seiler" birthdate="2012-07-15" gender="M" nation="SUI" swrid="5538025" athleteid="14221">
              <RESULTS>
                <RESULT eventid="1081" points="66" swimtime="00:01:59.25" resultid="14222" heatid="14561" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.87" />
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                    <SPLIT distance="75" swimtime="00:01:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="53" swimtime="00:02:26.50" resultid="14223" heatid="14616" lane="3" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.04" />
                    <SPLIT distance="50" swimtime="00:01:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="97" swimtime="00:01:37.55" resultid="14224" heatid="14668" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.03" />
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Dietiker" birthdate="2013-12-30" gender="M" nation="SUI" license="34378" swrid="5481964" athleteid="14042">
              <RESULTS>
                <RESULT eventid="1076" points="63" swimtime="00:00:55.77" resultid="14043" heatid="14536" lane="1" entrytime="00:01:00.81">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="206 - Unterwasserphase: Mehr als ein Delphinbeinschlag (Start) (Zeit: 12:00)" eventid="1090" status="DSQ" swimtime="00:01:04.24" resultid="14044" heatid="14591" lane="3" entrytime="00:01:30.16">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="58" swimtime="00:00:51.89" resultid="14045" heatid="14639" lane="4" entrytime="00:01:03.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mattea" lastname="Jakob" birthdate="2009-06-16" gender="F" nation="SUI" license="24839" swrid="5257621" athleteid="14107">
              <RESULTS>
                <RESULT eventid="1108" points="191" swimtime="00:01:34.79" resultid="14108" heatid="14686" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                    <SPLIT distance="75" swimtime="00:01:05.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="384" swimtime="00:01:15.48" resultid="14109" heatid="14714" lane="3" entrytime="00:01:13.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.98" />
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="75" swimtime="00:00:56.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="325" swimtime="00:01:30.62" resultid="14110" heatid="14744" lane="2" entrytime="00:01:30.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.13" />
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                    <SPLIT distance="75" swimtime="00:01:06.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="423" swimtime="00:01:06.93" resultid="14111" heatid="14774" lane="1" entrytime="00:01:09.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.79" />
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="75" swimtime="00:00:48.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessia" lastname="Fritschi" birthdate="2010-05-15" gender="F" nation="SUI" swrid="5168702" athleteid="14055">
              <RESULTS>
                <RESULT eventid="1078" points="160" swimtime="00:01:41.04" resultid="14056" heatid="14547" lane="1" entrytime="00:01:43.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.31" />
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                    <SPLIT distance="75" swimtime="00:01:16.35" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 12:18)" eventid="1092" status="DSQ" swimtime="00:01:55.33" resultid="14057" heatid="14604" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.92" />
                    <SPLIT distance="50" swimtime="00:00:53.71" />
                    <SPLIT distance="75" swimtime="00:01:24.72" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 14:13)" eventid="1102" status="DSQ" swimtime="00:01:21.20" resultid="14058" heatid="14657" lane="1" entrytime="00:01:22.72">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.92" />
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="75" swimtime="00:01:00.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lenja" lastname="Dietiker" birthdate="2013-03-11" gender="F" nation="SUI" swrid="5481965" athleteid="14046">
              <RESULTS>
                <RESULT eventid="1074" points="61" swimtime="00:01:05.00" resultid="14047" heatid="14527" lane="3" entrytime="00:01:19.00" />
                <RESULT eventid="1088" points="82" swimtime="00:01:05.49" resultid="14048" heatid="14586" lane="2" entrytime="00:01:10.30" />
                <RESULT eventid="1098" points="70" swimtime="00:00:55.50" resultid="14049" heatid="14633" lane="1" entrytime="00:01:01.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robin" lastname="Affentranger" birthdate="2004-03-19" gender="M" nation="SUI" license="24881" swrid="4745319" athleteid="13993">
              <RESULTS>
                <RESULT eventid="1111" points="511" swimtime="00:00:59.76" resultid="13994" heatid="14701" lane="1" entrytime="00:00:57.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                    <SPLIT distance="75" swimtime="00:00:43.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="599" swimtime="00:00:57.31" resultid="13995" heatid="14729" lane="2" entrytime="00:00:56.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.65" />
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                    <SPLIT distance="75" swimtime="00:00:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="544" swimtime="00:01:07.75" resultid="13996" heatid="14763" lane="4" entrytime="00:01:07.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.24" />
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                    <SPLIT distance="75" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="559" swimtime="00:00:54.53" resultid="13997" heatid="14797" lane="4" entrytime="00:00:53.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.80" />
                    <SPLIT distance="50" swimtime="00:00:26.54" />
                    <SPLIT distance="75" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="547" swimtime="00:00:27.16" resultid="14854" heatid="14802" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6683" points="507" swimtime="00:00:31.65" resultid="14866" heatid="14804" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6639" points="521" swimtime="00:00:27.03" resultid="14874" heatid="14806" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessia" lastname="Suter" birthdate="2012-08-23" gender="F" nation="SUI" license="25113" swrid="5439385" athleteid="14244">
              <RESULTS>
                <RESULT eventid="1078" points="118" swimtime="00:01:51.72" resultid="14245" heatid="14541" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.88" />
                    <SPLIT distance="50" swimtime="00:00:54.05" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Zeit: 12:14)" eventid="1092" status="DSQ" swimtime="00:02:06.00" resultid="14246" heatid="14595" lane="2" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.83" />
                    <SPLIT distance="75" swimtime="00:01:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="82" swimtime="00:01:55.28" resultid="14247" heatid="14647" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.05" />
                    <SPLIT distance="50" swimtime="00:01:00.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Campbell" birthdate="2010-10-24" gender="F" nation="SUI" license="25077" swrid="5351746" athleteid="14032">
              <RESULTS>
                <RESULT eventid="1068" points="255" swimtime="00:01:26.10" resultid="14033" heatid="14521" lane="3" entrytime="00:01:26.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.99" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:01:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="337" swimtime="00:01:18.84" resultid="14034" heatid="14553" lane="2" entrytime="00:01:20.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.63" />
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                    <SPLIT distance="75" swimtime="00:00:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="251" swimtime="00:01:38.77" resultid="14035" heatid="14607" lane="3" entrytime="00:01:39.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.72" />
                    <SPLIT distance="50" swimtime="00:00:47.23" />
                    <SPLIT distance="75" swimtime="00:01:13.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="322" swimtime="00:01:13.29" resultid="14036" heatid="14659" lane="1" entrytime="00:01:14.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.19" />
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yahya" lastname="Hussain" birthdate="2011-03-28" gender="M" nation="SUI" license="25087" swrid="5411013" athleteid="14097">
              <RESULTS>
                <RESULT eventid="1071" points="86" swimtime="00:01:48.00" resultid="14098" heatid="14523" lane="2" entrytime="00:02:15.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.71" />
                    <SPLIT distance="50" swimtime="00:00:50.04" />
                    <SPLIT distance="75" swimtime="00:01:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="173" swimtime="00:01:26.65" resultid="14099" heatid="14572" lane="1" entrytime="00:01:30.25">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.53" />
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="75" swimtime="00:01:06.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="113" swimtime="00:01:54.40" resultid="14100" heatid="14619" lane="3" entrytime="00:02:06.54">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.61" />
                    <SPLIT distance="50" swimtime="00:00:57.11" />
                    <SPLIT distance="75" swimtime="00:01:27.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="207" swimtime="00:01:15.97" resultid="14101" heatid="14679" lane="2" entrytime="00:01:17.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.09" />
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="75" swimtime="00:00:57.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roland" lastname="Neuenschwander" birthdate="2014-08-12" gender="M" nation="SUI" swrid="5551357" athleteid="14156">
              <RESULTS>
                <RESULT eventid="1076" points="57" swimtime="00:00:57.43" resultid="14157" heatid="14534" lane="3" entrytime="00:01:11.23">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="73" swimtime="00:01:00.30" resultid="14158" heatid="14593" lane="4" entrytime="00:01:07.09" />
                <RESULT eventid="1100" points="54" swimtime="00:00:53.06" resultid="14159" heatid="14639" lane="1" entrytime="00:00:56.39">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Radam" birthdate="2008-07-06" gender="M" nation="GER" license="24774" swrid="5185406" athleteid="14187">
              <RESULTS>
                <RESULT eventid="1111" points="377" swimtime="00:01:06.14" resultid="14188" heatid="14699" lane="1" entrytime="00:01:06.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.71" />
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="75" swimtime="00:00:47.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="396" swimtime="00:01:05.77" resultid="14189" heatid="14728" lane="3" entrytime="00:01:05.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.88" />
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="75" swimtime="00:00:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="345" swimtime="00:01:18.88" resultid="14190" heatid="14761" lane="2" entrytime="00:01:15.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.05" />
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="75" swimtime="00:00:57.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="407" swimtime="00:01:00.62" resultid="14191" heatid="14791" lane="2" entrytime="00:01:02.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.57" />
                    <SPLIT distance="50" swimtime="00:00:28.66" />
                    <SPLIT distance="75" swimtime="00:00:44.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Meta" lastname="Zimmermann" birthdate="2006-11-12" gender="F" nation="SUI" license="24843" swrid="5133832" athleteid="14280">
              <RESULTS>
                <RESULT eventid="1124" points="393" swimtime="00:01:25.08" resultid="14281" heatid="14748" lane="4" entrytime="00:01:24.45">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="75" swimtime="00:01:02.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="395" swimtime="00:01:08.45" resultid="14282" heatid="14779" lane="4" entrytime="00:01:03.61">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.09" />
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="75" swimtime="00:00:50.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Soyala" lastname="Déverin" birthdate="2007-10-01" gender="F" nation="SUI" license="25089" swrid="5382273" athleteid="14037">
              <RESULTS>
                <RESULT eventid="1108" points="418" swimtime="00:01:12.99" resultid="14038" heatid="14691" lane="4" entrytime="00:01:13.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="75" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="466" swimtime="00:01:10.76" resultid="14039" heatid="14715" lane="1" entrytime="00:01:11.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.06" />
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="75" swimtime="00:00:52.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="390" swimtime="00:01:25.29" resultid="14040" heatid="14748" lane="3" entrytime="00:01:23.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.02" />
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="75" swimtime="00:01:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="487" swimtime="00:01:03.86" resultid="14041" heatid="14778" lane="3" entrytime="00:01:04.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                    <SPLIT distance="75" swimtime="00:00:47.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lielle" lastname="Jakob" birthdate="2011-06-27" gender="F" nation="SUI" license="25079" swrid="5353514" athleteid="14102">
              <RESULTS>
                <RESULT eventid="1068" status="WDR" swimtime="00:00:00.00" resultid="14103" entrytime="00:02:00.00" />
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="14104" entrytime="00:01:46.74" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="14105" entrytime="00:01:55.80" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="14106" entrytime="00:01:31.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samantha" lastname="Stucki" birthdate="2010-04-20" gender="F" nation="SUI" license="29572" swrid="5451775" athleteid="14239">
              <RESULTS>
                <RESULT eventid="1068" points="309" swimtime="00:01:20.72" resultid="14240" heatid="14521" lane="1" entrytime="00:01:28.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.11" />
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="75" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="340" swimtime="00:01:18.58" resultid="14241" heatid="14553" lane="1" entrytime="00:01:21.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:59.53" />
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="251" swimtime="00:01:38.82" resultid="14242" heatid="14606" lane="2" entrytime="00:01:42.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.58" />
                    <SPLIT distance="50" swimtime="00:00:47.91" />
                    <SPLIT distance="75" swimtime="00:01:13.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="415" swimtime="00:01:07.32" resultid="14243" heatid="14661" lane="2" entrytime="00:01:07.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.27" />
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="75" swimtime="00:00:49.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Meier" birthdate="2008-07-06" gender="F" nation="SUI" license="24789" swrid="5257628" athleteid="14136">
              <RESULTS>
                <RESULT eventid="1114" points="315" swimtime="00:01:20.64" resultid="14137" heatid="14708" lane="1" entrytime="00:01:25.05">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.48" />
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="381" swimtime="00:01:09.31" resultid="14138" heatid="14771" lane="2" entrytime="00:01:11.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Vismara" birthdate="2005-10-04" gender="F" nation="ITA" license="24727" swrid="4964858" athleteid="14266">
              <RESULTS>
                <RESULT eventid="1108" points="737" swimtime="00:01:00.44" resultid="14267" heatid="14692" lane="2" entrytime="00:01:00.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.78" />
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="75" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="609" swimtime="00:01:04.75" resultid="14268" heatid="14716" lane="2" entrytime="00:01:01.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.02" />
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="75" swimtime="00:00:47.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="600" swimtime="00:01:13.93" resultid="14269" heatid="14750" lane="2" entrytime="00:01:14.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.81" />
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="75" swimtime="00:00:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="649" swimtime="00:00:58.03" resultid="14270" heatid="14781" lane="3" entrytime="00:00:58.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.13" />
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="75" swimtime="00:00:43.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="608" swimtime="00:00:30.21" resultid="14845" heatid="14801" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6681" points="566" swimtime="00:00:34.51" resultid="14862" heatid="14803" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6635" points="607" swimtime="00:00:28.79" resultid="14870" heatid="14805" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6637" points="653" swimtime="00:00:26.43" resultid="14876" heatid="14807" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manon" lastname="Bircher" birthdate="2011-04-24" gender="F" nation="SUI" license="29355" swrid="5456692" athleteid="14022">
              <RESULTS>
                <RESULT eventid="1068" points="143" swimtime="00:01:44.24" resultid="14023" heatid="14519" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.41" />
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                    <SPLIT distance="75" swimtime="00:01:13.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="227" swimtime="00:01:29.97" resultid="14024" heatid="14550" lane="2" entrytime="00:01:35.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.16" />
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="75" swimtime="00:01:07.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="270" swimtime="00:01:36.38" resultid="14025" heatid="14607" lane="4" entrytime="00:01:41.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.86" />
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="75" swimtime="00:01:11.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="281" swimtime="00:01:16.67" resultid="14026" heatid="14657" lane="2" entrytime="00:01:22.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="75" swimtime="00:00:56.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mila" lastname="Binder" birthdate="2012-07-14" gender="F" nation="SUI" swrid="5449263" athleteid="14018">
              <RESULTS>
                <RESULT eventid="1078" points="114" swimtime="00:01:52.88" resultid="14019" heatid="14541" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.62" />
                    <SPLIT distance="75" swimtime="00:01:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="134" swimtime="00:02:01.80" resultid="14020" heatid="14597" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.46" />
                    <SPLIT distance="50" swimtime="00:00:55.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="118" swimtime="00:01:42.41" resultid="14021" heatid="14646" lane="4" entrytime="00:01:56.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.54" />
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="75" swimtime="00:01:15.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Moira" lastname="Gämperle" birthdate="2011-01-21" gender="F" nation="SUI" license="25120" swrid="5439383" athleteid="14059">
              <RESULTS>
                <RESULT eventid="1068" points="137" swimtime="00:01:45.88" resultid="14060" heatid="14520" lane="1" entrytime="00:01:40.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.59" />
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="75" swimtime="00:01:15.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="222" swimtime="00:01:30.58" resultid="14061" heatid="14551" lane="3" entrytime="00:01:35.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.71" />
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="75" swimtime="00:01:07.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="156" swimtime="00:01:55.62" resultid="14062" heatid="14602" lane="1" entrytime="00:01:56.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.72" />
                    <SPLIT distance="50" swimtime="00:00:53.81" />
                    <SPLIT distance="75" swimtime="00:01:25.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="226" swimtime="00:01:22.39" resultid="14063" heatid="14657" lane="4" entrytime="00:01:22.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                    <SPLIT distance="75" swimtime="00:01:01.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Radam" birthdate="2004-06-06" gender="M" nation="SUI" license="24760" swrid="4830858" athleteid="14182">
              <RESULTS>
                <RESULT eventid="1111" points="552" swimtime="00:00:58.24" resultid="14183" heatid="14701" lane="2" entrytime="00:00:56.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.59" />
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                    <SPLIT distance="75" swimtime="00:00:43.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="612" swimtime="00:00:56.92" resultid="14184" heatid="14729" lane="3" entrytime="00:00:56.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.52" />
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                    <SPLIT distance="75" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="466" swimtime="00:01:11.36" resultid="14185" heatid="14755" lane="2" entrytime="00:01:35.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="75" swimtime="00:00:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="562" swimtime="00:00:54.43" resultid="14186" heatid="14797" lane="1" entrytime="00:00:52.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.40" />
                    <SPLIT distance="50" swimtime="00:00:26.53" />
                    <SPLIT distance="75" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="542" swimtime="00:00:27.25" resultid="14857" heatid="14843" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6683" points="495" swimtime="00:00:31.91" resultid="14869" heatid="14804" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6639" points="560" swimtime="00:00:26.38" resultid="14875" heatid="14806" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6679" points="564" swimtime="00:00:24.39" resultid="14879" heatid="14808" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="527" swimtime="00:01:51.91" resultid="14283" heatid="14736" lane="2" entrytime="00:01:47.83">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.43" />
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                    <SPLIT distance="75" swimtime="00:00:41.49" />
                    <SPLIT distance="100" swimtime="00:00:58.87" />
                    <SPLIT distance="125" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:25.27" />
                    <SPLIT distance="175" swimtime="00:01:38.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13993" number="1" />
                    <RELAYPOSITION athleteid="14197" number="2" />
                    <RELAYPOSITION athleteid="14182" number="3" />
                    <RELAYPOSITION athleteid="14252" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="205" swimtime="00:02:18.59" resultid="14813" heatid="14818" lane="3" entrytime="00:02:15.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:08.39" />
                    <SPLIT distance="125" swimtime="00:01:26.07" />
                    <SPLIT distance="150" swimtime="00:01:45.44" />
                    <SPLIT distance="175" swimtime="00:02:01.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14163" number="1" />
                    <RELAYPOSITION athleteid="14097" number="2" />
                    <RELAYPOSITION athleteid="14050" number="3" />
                    <RELAYPOSITION athleteid="14168" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1122" points="429" swimtime="00:01:59.91" resultid="14284" heatid="14735" lane="1" entrytime="00:02:26.68">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.34" />
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="75" swimtime="00:00:44.89" />
                    <SPLIT distance="100" swimtime="00:01:02.48" />
                    <SPLIT distance="125" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:01:32.35" />
                    <SPLIT distance="175" swimtime="00:01:45.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14187" number="1" />
                    <RELAYPOSITION athleteid="13988" number="2" />
                    <RELAYPOSITION athleteid="14173" number="3" />
                    <RELAYPOSITION athleteid="14261" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1086" points="161" swimtime="00:02:30.35" resultid="14814" heatid="14583" lane="3" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="75" swimtime="00:00:58.41" />
                    <SPLIT distance="100" swimtime="00:01:17.17" />
                    <SPLIT distance="125" swimtime="00:01:35.18" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                    <SPLIT distance="175" swimtime="00:02:12.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14064" number="1" />
                    <RELAYPOSITION athleteid="14116" number="2" />
                    <RELAYPOSITION athleteid="14178" number="3" />
                    <RELAYPOSITION athleteid="14027" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1086" points="91" swimtime="00:03:01.56" resultid="14815" heatid="14582" lane="4" entrytime="00:02:56.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.36" />
                    <SPLIT distance="50" swimtime="00:00:51.86" />
                    <SPLIT distance="75" swimtime="00:01:12.70" />
                    <SPLIT distance="100" swimtime="00:01:34.26" />
                    <SPLIT distance="125" swimtime="00:01:55.16" />
                    <SPLIT distance="150" swimtime="00:02:18.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14068" number="1" />
                    <RELAYPOSITION athleteid="14221" number="2" />
                    <RELAYPOSITION athleteid="14081" number="3" />
                    <RELAYPOSITION athleteid="14093" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1086" points="66" swimtime="00:03:21.69" resultid="14816" heatid="14581" lane="3" entrytime="00:03:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.44" />
                    <SPLIT distance="75" swimtime="00:01:14.47" />
                    <SPLIT distance="100" swimtime="00:01:43.41" />
                    <SPLIT distance="125" swimtime="00:02:06.21" />
                    <SPLIT distance="150" swimtime="00:02:32.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14125" number="1" />
                    <RELAYPOSITION athleteid="14156" number="2" />
                    <RELAYPOSITION athleteid="14152" number="3" />
                    <RELAYPOSITION athleteid="14042" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="584" swimtime="00:02:02.47" resultid="14285" heatid="14733" lane="2" entrytime="00:02:00.71">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="75" swimtime="00:00:46.32" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="125" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:01:35.38" />
                    <SPLIT distance="175" swimtime="00:01:48.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14275" number="1" />
                    <RELAYPOSITION athleteid="14266" number="2" />
                    <RELAYPOSITION athleteid="14192" number="3" />
                    <RELAYPOSITION athleteid="14003" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="342" swimtime="00:02:12.25" resultid="14809" heatid="14817" lane="2" entrytime="00:02:09.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.55" />
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="75" swimtime="00:00:47.05" />
                    <SPLIT distance="100" swimtime="00:01:06.05" />
                    <SPLIT distance="125" swimtime="00:01:22.10" />
                    <SPLIT distance="150" swimtime="00:01:40.32" />
                    <SPLIT distance="175" swimtime="00:01:55.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14239" number="1" />
                    <RELAYPOSITION athleteid="14212" number="2" />
                    <RELAYPOSITION athleteid="14022" number="3" />
                    <RELAYPOSITION athleteid="14032" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer ...), Schwimmer 3" eventid="1120" status="DSQ" swimtime="00:02:10.59" resultid="14286" heatid="14733" lane="3" entrytime="00:02:10.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.78" />
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="75" swimtime="00:00:52.24" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="125" swimtime="00:01:25.78" />
                    <SPLIT distance="150" swimtime="00:01:42.88" />
                    <SPLIT distance="175" swimtime="00:01:56.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14139" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="14008" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="14037" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="14076" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1084" points="186" swimtime="00:02:41.99" resultid="14810" heatid="14580" lane="2" entrytime="00:02:27.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.31" />
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                    <SPLIT distance="75" swimtime="00:01:00.27" />
                    <SPLIT distance="100" swimtime="00:01:26.58" />
                    <SPLIT distance="125" swimtime="00:01:43.92" />
                    <SPLIT distance="150" swimtime="00:02:03.15" />
                    <SPLIT distance="175" swimtime="00:02:21.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14120" number="1" />
                    <RELAYPOSITION athleteid="14234" number="2" />
                    <RELAYPOSITION athleteid="14055" number="3" />
                    <RELAYPOSITION athleteid="14059" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1120" points="329" swimtime="00:02:28.17" resultid="14287" heatid="14732" lane="1" entrytime="00:02:26.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="75" swimtime="00:00:58.94" />
                    <SPLIT distance="100" swimtime="00:01:21.91" />
                    <SPLIT distance="125" swimtime="00:01:38.38" />
                    <SPLIT distance="150" swimtime="00:01:57.84" />
                    <SPLIT distance="175" swimtime="00:02:12.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14011" number="1" />
                    <RELAYPOSITION athleteid="14136" number="2" />
                    <RELAYPOSITION athleteid="14229" number="3" />
                    <RELAYPOSITION athleteid="14107" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1084" points="94" swimtime="00:03:22.80" resultid="14811" heatid="14577" lane="1" entrytime="00:03:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.38" />
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="75" swimtime="00:01:13.76" />
                    <SPLIT distance="100" swimtime="00:01:41.43" />
                    <SPLIT distance="125" swimtime="00:02:07.98" />
                    <SPLIT distance="150" swimtime="00:02:38.57" />
                    <SPLIT distance="175" swimtime="00:03:00.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14244" number="1" />
                    <RELAYPOSITION athleteid="14132" number="2" />
                    <RELAYPOSITION athleteid="14014" number="3" />
                    <RELAYPOSITION athleteid="14018" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="4">
              <RESULTS>
                <RESULT eventid="1084" points="44" swimtime="00:04:20.77" resultid="14812" heatid="14576" lane="3" entrytime="00:03:52.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.99" />
                    <SPLIT distance="50" swimtime="00:00:55.51" />
                    <SPLIT distance="75" swimtime="00:01:24.44" />
                    <SPLIT distance="100" swimtime="00:02:01.82" />
                    <SPLIT distance="125" swimtime="00:02:40.40" />
                    <SPLIT distance="150" swimtime="00:03:22.82" />
                    <SPLIT distance="175" swimtime="00:03:49.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14046" number="1" />
                    <RELAYPOSITION athleteid="14271" number="2" />
                    <RELAYPOSITION athleteid="14148" number="3" />
                    <RELAYPOSITION athleteid="14225" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="OW88" nation="SUI" region="RSR" clubid="12486" swrid="65577" name="Schwimmverein Oberwallis" shortname="ow88">
          <ATHLETES>
            <ATHLETE firstname="Milena" lastname="Lengen" birthdate="2006-07-11" gender="F" nation="SUI" license="24396" swrid="5222669" athleteid="12516">
              <RESULTS>
                <RESULT eventid="1108" points="253" swimtime="00:01:26.27" resultid="12517" heatid="14686" lane="1" entrytime="00:01:30.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.35" />
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="75" swimtime="00:01:01.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="349" swimtime="00:01:28.49" resultid="12518" heatid="14747" lane="4" entrytime="00:01:26.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.94" />
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                    <SPLIT distance="75" swimtime="00:01:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="344" swimtime="00:01:11.66" resultid="12519" heatid="14772" lane="2" entrytime="00:01:11.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.84" />
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="75" swimtime="00:00:53.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Silas" lastname="Stump" birthdate="2010-11-06" gender="M" nation="SUI" license="24536" swrid="5479918" athleteid="12557">
              <RESULTS>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...) (Zeit: 9:10)" eventid="1071" status="DSQ" swimtime="00:02:06.77" resultid="12558" heatid="14524" lane="1" entrytime="00:02:11.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.59" />
                    <SPLIT distance="50" swimtime="00:00:56.71" />
                    <SPLIT distance="75" swimtime="00:01:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="114" swimtime="00:01:39.46" resultid="12559" heatid="14565" lane="2" entrytime="00:01:49.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.86" />
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="206 - Unterwasserphase: Mehr als ein Delphinbeinschlag (Start) (Zeit: 13:10)" eventid="1095" status="DSQ" swimtime="00:01:55.25" resultid="12560" heatid="14623" lane="4" entrytime="00:01:53.59">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.28" />
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                    <SPLIT distance="75" swimtime="00:01:24.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="104" swimtime="00:01:35.29" resultid="12561" heatid="14676" lane="4" entrytime="00:01:30.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.71" />
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Slatincic" birthdate="2012-08-06" gender="F" nation="SUI" license="24274" swrid="5529905" athleteid="12530">
              <RESULTS>
                <RESULT eventid="1078" points="119" swimtime="00:01:51.57" resultid="12531" heatid="14540" lane="1" entrytime="00:02:05.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.54" />
                    <SPLIT distance="50" swimtime="00:00:54.86" />
                    <SPLIT distance="75" swimtime="00:01:25.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="100" swimtime="00:02:13.91" resultid="12532" heatid="14596" lane="2" entrytime="00:02:20.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.13" />
                    <SPLIT distance="50" swimtime="00:01:02.62" />
                    <SPLIT distance="75" swimtime="00:01:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="117" swimtime="00:01:42.69" resultid="12533" heatid="14650" lane="4" entrytime="00:01:38.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.31" />
                    <SPLIT distance="50" swimtime="00:00:48.38" />
                    <SPLIT distance="75" swimtime="00:01:16.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Jäger" birthdate="2012-11-03" gender="F" nation="SUI" license="24216" swrid="5529894" athleteid="12508">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 9:57)" eventid="1078" status="DSQ" swimtime="00:02:25.12" resultid="12509" heatid="14538" lane="2" entrytime="00:02:23.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.34" />
                    <SPLIT distance="50" swimtime="00:01:09.21" />
                    <SPLIT distance="75" swimtime="00:01:47.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="97" swimtime="00:02:15.50" resultid="12510" heatid="14595" lane="4" entrytime="00:02:40.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.02" />
                    <SPLIT distance="50" swimtime="00:01:02.59" />
                    <SPLIT distance="75" swimtime="00:01:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="42" swimtime="00:02:24.55" resultid="12511" heatid="14643" lane="1" entrytime="00:02:22.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.65" />
                    <SPLIT distance="50" swimtime="00:01:01.78" />
                    <SPLIT distance="75" swimtime="00:01:44.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Jossen" birthdate="2007-08-31" gender="F" nation="SUI" license="35874" swrid="5486806" athleteid="12512">
              <RESULTS>
                <RESULT eventid="1114" points="165" swimtime="00:01:39.92" resultid="12513" heatid="14705" lane="4" entrytime="00:01:35.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.51" />
                    <SPLIT distance="50" swimtime="00:00:47.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="208" swimtime="00:01:45.10" resultid="12514" heatid="14740" lane="4" entrytime="00:01:48.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.65" />
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                    <SPLIT distance="75" swimtime="00:01:16.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="171" swimtime="00:01:30.41" resultid="12515" heatid="14766" lane="2" entrytime="00:01:26.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.03" />
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="75" swimtime="00:01:06.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ilaria" lastname="Battaglia" birthdate="2011-12-18" gender="F" nation="SUI" athleteid="12487">
              <RESULTS>
                <RESULT comment="204 - Starten vor dem Startkommando" eventid="1078" status="DSQ" swimtime="00:02:18.94" resultid="12488" heatid="14538" lane="1" entrytime="00:02:29.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.50" />
                    <SPLIT distance="50" swimtime="00:01:04.12" />
                    <SPLIT distance="75" swimtime="00:01:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="65" swimtime="00:02:34.57" resultid="12489" heatid="14595" lane="1" entrytime="00:02:38.08">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.40" />
                    <SPLIT distance="50" swimtime="00:01:10.61" />
                    <SPLIT distance="75" swimtime="00:01:53.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="79" swimtime="00:01:56.68" resultid="12490" heatid="14644" lane="1" entrytime="00:02:11.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.66" />
                    <SPLIT distance="50" swimtime="00:00:54.92" />
                    <SPLIT distance="75" swimtime="00:01:27.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ladina" lastname="Stoffel" birthdate="2010-08-13" gender="F" nation="SUI" license="24116" swrid="5336558" athleteid="12544">
              <RESULTS>
                <RESULT eventid="1068" points="155" swimtime="00:01:41.52" resultid="12545" heatid="14517" lane="1" entrytime="00:02:09.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.42" />
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                    <SPLIT distance="75" swimtime="00:01:14.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="212" swimtime="00:01:32.04" resultid="12546" heatid="14544" lane="2" entrytime="00:01:46.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.31" />
                    <SPLIT distance="75" swimtime="00:01:09.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="272" swimtime="00:01:36.20" resultid="12547" heatid="14606" lane="1" entrytime="00:01:42.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.90" />
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                    <SPLIT distance="75" swimtime="00:01:10.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="212" swimtime="00:01:24.19" resultid="12548" heatid="14652" lane="2" entrytime="00:01:28.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.39" />
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="75" swimtime="00:01:02.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elio" lastname="Vogel" birthdate="2009-10-07" gender="M" nation="SUI" license="24126" swrid="4590434" athleteid="12562">
              <RESULTS>
                <RESULT eventid="1111" points="81" swimtime="00:01:50.12" resultid="12563" heatid="14695" lane="1" entrytime="00:01:55.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.77" />
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                    <SPLIT distance="75" swimtime="00:01:23.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="131" swimtime="00:01:34.96" resultid="12564" heatid="14719" lane="2" entrytime="00:01:38.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.49" />
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="121" swimtime="00:01:51.84" resultid="12565" heatid="14753" lane="1" entrytime="00:01:55.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.38" />
                    <SPLIT distance="50" swimtime="00:00:53.68" />
                    <SPLIT distance="75" swimtime="00:01:22.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="116" swimtime="00:01:32.10" resultid="12566" heatid="14784" lane="3" entrytime="00:01:29.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.86" />
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Walker" birthdate="2011-01-10" gender="M" nation="SUI" license="24440" swrid="5418201" athleteid="12567">
              <RESULTS>
                <RESULT eventid="1071" points="70" swimtime="00:01:55.92" resultid="12568" heatid="14524" lane="2" entrytime="00:01:53.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.99" />
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                    <SPLIT distance="75" swimtime="00:01:25.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="404 - Nicht in Rückenlage angeschlagen (Ziel) (Zeit: 10:46)" eventid="1081" status="DSQ" swimtime="00:01:38.26" resultid="12569" heatid="14570" lane="1" entrytime="00:01:37.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="151" swimtime="00:01:43.86" resultid="12570" heatid="14626" lane="2" entrytime="00:01:44.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.19" />
                    <SPLIT distance="50" swimtime="00:00:49.44" />
                    <SPLIT distance="75" swimtime="00:01:17.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="136" swimtime="00:01:27.30" resultid="12571" heatid="14677" lane="4" entrytime="00:01:28.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.68" />
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="75" swimtime="00:01:04.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Stoffel" birthdate="2012-10-12" gender="M" nation="SUI" license="24677" swrid="5531321" athleteid="12549">
              <RESULTS>
                <RESULT eventid="1081" points="45" swimtime="00:02:15.22" resultid="12550" heatid="14559" lane="4" entrytime="00:02:32.62">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.36" />
                    <SPLIT distance="50" swimtime="00:01:04.11" />
                    <SPLIT distance="75" swimtime="00:01:42.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="62" swimtime="00:02:19.17" resultid="12551" heatid="14614" lane="2" entrytime="00:02:40.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.76" />
                    <SPLIT distance="50" swimtime="00:01:08.10" />
                    <SPLIT distance="75" swimtime="00:01:43.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="41" swimtime="00:02:09.97" resultid="12552" heatid="14666" lane="3" entrytime="00:02:05.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.20" />
                    <SPLIT distance="50" swimtime="00:00:57.64" />
                    <SPLIT distance="75" swimtime="00:01:35.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lian" lastname="Stump" birthdate="2012-08-05" gender="M" nation="SUI" license="24279" swrid="5418189" athleteid="12553">
              <RESULTS>
                <RESULT eventid="1081" points="86" swimtime="00:01:49.09" resultid="12554" heatid="14563" lane="4" entrytime="00:02:01.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.59" />
                    <SPLIT distance="50" swimtime="00:00:53.08" />
                    <SPLIT distance="75" swimtime="00:01:22.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="91" swimtime="00:02:03.01" resultid="12555" heatid="14618" lane="3" entrytime="00:02:09.38">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.47" />
                    <SPLIT distance="50" swimtime="00:00:57.18" />
                    <SPLIT distance="75" swimtime="00:01:29.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="84" swimtime="00:01:42.37" resultid="12556" heatid="14672" lane="4" entrytime="00:01:37.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.19" />
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                    <SPLIT distance="75" swimtime="00:01:16.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Imboden" birthdate="2012-03-12" gender="F" nation="SUI" license="24207" swrid="5305724" athleteid="12504">
              <RESULTS>
                <RESULT eventid="1078" points="69" swimtime="00:02:13.42" resultid="12505" heatid="14539" lane="3" entrytime="00:02:10.38">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.81" />
                    <SPLIT distance="50" swimtime="00:01:02.47" />
                    <SPLIT distance="75" swimtime="00:01:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="113" swimtime="00:02:08.78" resultid="12506" heatid="14596" lane="3" entrytime="00:02:21.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.68" />
                    <SPLIT distance="50" swimtime="00:01:01.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="51" swimtime="00:02:14.92" resultid="12507" heatid="14643" lane="2" entrytime="00:02:12.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.00" />
                    <SPLIT distance="50" swimtime="00:00:59.97" />
                    <SPLIT distance="75" swimtime="00:01:37.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elias" lastname="Steffen" birthdate="2011-10-02" gender="M" nation="SUI" license="24427" swrid="5418192" athleteid="12534">
              <RESULTS>
                <RESULT eventid="1071" points="71" swimtime="00:01:55.28" resultid="12535" heatid="14523" lane="3" entrytime="00:02:17.15">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.48" />
                    <SPLIT distance="50" swimtime="00:00:49.05" />
                    <SPLIT distance="75" swimtime="00:01:21.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="114" swimtime="00:01:39.46" resultid="12536" heatid="14566" lane="2" entrytime="00:01:48.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.86" />
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="121" swimtime="00:01:51.58" resultid="12537" heatid="14624" lane="1" entrytime="00:01:52.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.32" />
                    <SPLIT distance="50" swimtime="00:00:53.71" />
                    <SPLIT distance="75" swimtime="00:01:23.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="127" swimtime="00:01:29.32" resultid="12538" heatid="14672" lane="1" entrytime="00:01:36.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.82" />
                    <SPLIT distance="50" swimtime="00:01:29.95" />
                    <SPLIT distance="75" swimtime="00:01:08.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Mengis" birthdate="2007-09-10" gender="F" nation="SUI" license="24404" swrid="5222672" athleteid="12525">
              <RESULTS>
                <RESULT eventid="1108" points="296" swimtime="00:01:21.88" resultid="12526" heatid="14688" lane="1" entrytime="00:01:22.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.12" />
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="75" swimtime="00:00:58.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="352" swimtime="00:01:17.68" resultid="12527" heatid="14713" lane="2" entrytime="00:01:14.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.73" />
                    <SPLIT distance="50" swimtime="00:00:36.62" />
                    <SPLIT distance="75" swimtime="00:00:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="254" swimtime="00:01:38.45" resultid="12528" heatid="14742" lane="4" entrytime="00:01:36.55">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.30" />
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                    <SPLIT distance="75" swimtime="00:01:12.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="407" swimtime="00:01:07.80" resultid="12529" heatid="14775" lane="1" entrytime="00:01:07.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.20" />
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="75" swimtime="00:00:50.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benedikt" lastname="Brigger" birthdate="2007-09-29" gender="M" nation="SUI" license="24341" swrid="5222670" athleteid="12495">
              <RESULTS>
                <RESULT eventid="1111" points="247" swimtime="00:01:16.13" resultid="12496" heatid="14696" lane="3" entrytime="00:01:25.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.89" />
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="75" swimtime="00:00:55.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="280" swimtime="00:01:24.51" resultid="12497" heatid="14758" lane="3" entrytime="00:01:27.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.84" />
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="75" swimtime="00:01:02.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="331" swimtime="00:01:04.91" resultid="12498" heatid="14790" lane="3" entrytime="00:01:04.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.83" />
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="75" swimtime="00:00:48.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessandra" lastname="Mangisch" birthdate="2009-09-05" gender="F" nation="SUI" license="24399" swrid="5348936" athleteid="12520">
              <RESULTS>
                <RESULT eventid="1108" points="172" swimtime="00:01:38.12" resultid="12521" heatid="14685" lane="4" entrytime="00:01:36.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.89" />
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                    <SPLIT distance="75" swimtime="00:01:10.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="247" swimtime="00:01:27.37" resultid="12522" heatid="14705" lane="2" entrytime="00:01:32.67">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.01" />
                    <SPLIT distance="50" swimtime="00:00:42.27" />
                    <SPLIT distance="75" swimtime="00:01:05.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="263" swimtime="00:01:37.33" resultid="12523" heatid="14741" lane="4" entrytime="00:01:39.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.70" />
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="75" swimtime="00:01:13.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="263" swimtime="00:01:18.38" resultid="12524" heatid="14769" lane="4" entrytime="00:01:17.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.75" />
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="75" swimtime="00:00:58.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Neele" lastname="Heinen" birthdate="2011-06-15" gender="F" nation="SUI" license="24585" swrid="5418199" athleteid="12499">
              <RESULTS>
                <RESULT eventid="1068" points="141" swimtime="00:01:44.77" resultid="12500" heatid="14519" lane="1" entrytime="00:01:45.37">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.95" />
                    <SPLIT distance="50" swimtime="00:00:48.97" />
                    <SPLIT distance="75" swimtime="00:01:18.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="188" swimtime="00:01:35.78" resultid="12501" heatid="14547" lane="4" entrytime="00:01:44.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.61" />
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="75" swimtime="00:01:11.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="188" swimtime="00:01:48.78" resultid="12502" heatid="14597" lane="3" entrytime="00:02:11.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.21" />
                    <SPLIT distance="50" swimtime="00:00:51.82" />
                    <SPLIT distance="75" swimtime="00:01:19.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="239" swimtime="00:01:20.95" resultid="12503" heatid="14654" lane="3" entrytime="00:01:26.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.05" />
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="75" swimtime="00:01:00.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Steffen" birthdate="2014-01-11" gender="F" nation="SUI" license="24276" swrid="5310814" athleteid="12539">
              <RESULTS>
                <RESULT eventid="1064" points="49" swimtime="00:01:06.55" resultid="14819" heatid="14514" lane="3" entrytime="00:00:59.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="104" swimtime="00:00:54.32" resultid="14820" heatid="14532" lane="4" entrytime="00:00:54.80" />
                <RESULT eventid="1088" points="117" swimtime="00:00:58.37" resultid="14821" heatid="14587" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="117" swimtime="00:00:46.77" resultid="14822" heatid="14635" lane="2" entrytime="00:00:50.06">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Walker" birthdate="2010-12-26" gender="F" nation="SUI" license="38143" swrid="5529907" athleteid="12572">
              <RESULTS>
                <RESULT eventid="1068" points="151" swimtime="00:01:42.54" resultid="12573" heatid="14517" lane="2" entrytime="00:01:59.18" />
                <RESULT eventid="1078" points="218" swimtime="00:01:31.16" resultid="12574" heatid="14547" lane="3" entrytime="00:01:42.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:31.18" />
                    <SPLIT distance="75" swimtime="00:01:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="204" swimtime="00:01:45.84" resultid="12575" heatid="14601" lane="4" entrytime="00:02:00.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.93" />
                    <SPLIT distance="50" swimtime="00:00:50.91" />
                    <SPLIT distance="75" swimtime="00:01:18.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="234" swimtime="00:01:21.46" resultid="12576" heatid="14651" lane="1" entrytime="00:01:35.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.78" />
                    <SPLIT distance="50" swimtime="00:00:39.46" />
                    <SPLIT distance="75" swimtime="00:01:00.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Bregy" birthdate="2008-12-08" gender="F" nation="SUI" license="35151" swrid="5486795" athleteid="12491">
              <RESULTS>
                <RESULT eventid="1108" points="85" swimtime="00:02:03.86" resultid="12492" heatid="14684" lane="1" entrytime="00:01:50.09">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.98" />
                    <SPLIT distance="50" swimtime="00:00:54.89" />
                    <SPLIT distance="75" swimtime="00:01:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="250" swimtime="00:01:38.89" resultid="12493" heatid="14740" lane="1" entrytime="00:01:42.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.68" />
                    <SPLIT distance="50" swimtime="00:00:47.68" />
                    <SPLIT distance="75" swimtime="00:01:13.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="209" swimtime="00:01:24.60" resultid="12494" heatid="14767" lane="2" entrytime="00:01:22.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.88" />
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="75" swimtime="00:01:03.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="117" swimtime="00:02:46.96" resultid="12577" heatid="14582" lane="3" entrytime="00:02:45.18">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.86" />
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="75" swimtime="00:01:03.68" />
                    <SPLIT distance="100" swimtime="00:01:27.94" />
                    <SPLIT distance="125" swimtime="00:01:46.92" />
                    <SPLIT distance="150" swimtime="00:02:07.93" />
                    <SPLIT distance="175" swimtime="00:02:26.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12557" number="1" />
                    <RELAYPOSITION athleteid="12553" number="2" />
                    <RELAYPOSITION athleteid="12534" number="3" />
                    <RELAYPOSITION athleteid="12567" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="218" swimtime="00:02:33.67" resultid="12578" heatid="14578" lane="3" entrytime="00:02:49.73">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.03" />
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="75" swimtime="00:00:53.08" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="125" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:01:57.02" />
                    <SPLIT distance="175" swimtime="00:02:14.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12499" number="1" />
                    <RELAYPOSITION athleteid="12572" number="2" />
                    <RELAYPOSITION athleteid="12530" number="3" />
                    <RELAYPOSITION athleteid="12544" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="308" swimtime="00:02:31.45" resultid="12579" heatid="14731" lane="2" entrytime="00:02:33.97">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.27" />
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="75" swimtime="00:00:52.77" />
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                    <SPLIT distance="125" swimtime="00:01:32.10" />
                    <SPLIT distance="150" swimtime="00:01:54.73" />
                    <SPLIT distance="175" swimtime="00:02:12.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12525" number="1" />
                    <RELAYPOSITION athleteid="12516" number="2" />
                    <RELAYPOSITION athleteid="12520" number="3" />
                    <RELAYPOSITION athleteid="12491" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1084" points="74" swimtime="00:03:39.72" resultid="12580" heatid="14576" lane="1" entrytime="00:04:09.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.85" />
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                    <SPLIT distance="75" swimtime="00:01:16.68" />
                    <SPLIT distance="100" swimtime="00:01:52.28" />
                    <SPLIT distance="125" swimtime="00:03:08.76" />
                    <SPLIT distance="150" swimtime="00:02:44.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12539" number="1" />
                    <RELAYPOSITION athleteid="12508" number="2" />
                    <RELAYPOSITION athleteid="12487" number="3" />
                    <RELAYPOSITION athleteid="12504" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BIEL" nation="SUI" region="RZW" clubid="12682" swrid="65714" name="Swim Team Biel-Bienne" shortname="Biel">
          <ATHLETES>
            <ATHLETE firstname="Eléna" lastname="Zaffino" birthdate="2010-05-11" gender="F" nation="ITA" license="7147" swrid="5255766" athleteid="12812">
              <RESULTS>
                <RESULT eventid="1068" points="211" swimtime="00:01:31.71" resultid="12813" heatid="14522" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="316" swimtime="00:01:20.56" resultid="12814" heatid="14553" lane="3" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.16" />
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="75" swimtime="00:01:00.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="285" swimtime="00:01:34.74" resultid="12815" heatid="14608" lane="3" entrytime="00:01:36.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.94" />
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="75" swimtime="00:01:10.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="320" swimtime="00:01:13.46" resultid="12816" heatid="14659" lane="2" entrytime="00:01:13.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Dumitru" birthdate="2013-09-22" gender="M" nation="ROU" license="42543" athleteid="12692">
              <RESULTS>
                <RESULT eventid="1076" status="WDR" swimtime="00:00:00.00" resultid="12693" entrytime="00:00:56.63" entrycourse="SCM" />
                <RESULT eventid="1090" status="WDR" swimtime="00:00:00.00" resultid="12694" entrytime="00:01:10.00" />
                <RESULT eventid="1100" status="WDR" swimtime="00:00:00.00" resultid="12695" entrytime="00:00:53.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jaron" lastname="Schwab" birthdate="2011-01-24" gender="M" nation="SUI" license="7164" swrid="5335435" athleteid="12790">
              <RESULTS>
                <RESULT eventid="1071" points="111" swimtime="00:01:39.26" resultid="12791" heatid="14525" lane="2" entrytime="00:01:43.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.95" />
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                    <SPLIT distance="75" swimtime="00:01:10.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="142" swimtime="00:01:32.46" resultid="12792" heatid="14572" lane="4" entrytime="00:01:30.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.05" />
                    <SPLIT distance="50" swimtime="00:00:46.05" />
                    <SPLIT distance="75" swimtime="00:01:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="181" swimtime="00:01:37.66" resultid="12793" heatid="14628" lane="3" entrytime="00:01:37.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.56" />
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="75" swimtime="00:01:12.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="215" swimtime="00:01:14.96" resultid="12794" heatid="14679" lane="3" entrytime="00:01:18.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.96" />
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="75" swimtime="00:00:57.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livio" lastname="Milandri" birthdate="2011-09-29" gender="M" nation="FRA" license="7183" swrid="5411051" athleteid="12759">
              <RESULTS>
                <RESULT eventid="1081" points="102" swimtime="00:01:43.36" resultid="12760" heatid="14568" lane="1" entrytime="00:01:44.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.52" />
                    <SPLIT distance="50" swimtime="00:00:50.29" />
                    <SPLIT distance="75" swimtime="00:01:17.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="116" swimtime="00:01:53.40" resultid="12761" heatid="14622" lane="3" entrytime="00:01:54.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.06" />
                    <SPLIT distance="50" swimtime="00:00:53.36" />
                    <SPLIT distance="75" swimtime="00:01:23.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="103" swimtime="00:01:35.59" resultid="12762" heatid="14673" lane="4" entrytime="00:01:36.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.87" />
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                    <SPLIT distance="75" swimtime="00:01:10.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dimitri" lastname="König" birthdate="2011-12-15" gender="M" nation="SUI" license="7144" swrid="5411041" athleteid="12734">
              <RESULTS>
                <RESULT eventid="1081" points="98" swimtime="00:01:44.80" resultid="12735" heatid="14568" lane="4" entrytime="00:01:44.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.97" />
                    <SPLIT distance="50" swimtime="00:00:50.13" />
                    <SPLIT distance="75" swimtime="00:01:18.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="307 - Unterwasserphase: Mehr als ein Delphinbeinschlag (Wende 1) (Zeit: 13:11)" eventid="1095" status="DSQ" swimtime="00:01:48.75" resultid="12736" heatid="14624" lane="4" entrytime="00:01:52.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.73" />
                    <SPLIT distance="50" swimtime="00:00:52.32" />
                    <SPLIT distance="75" swimtime="00:01:20.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="104" swimtime="00:01:35.47" resultid="12737" heatid="14674" lane="2" entrytime="00:01:32.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.40" />
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="75" swimtime="00:01:10.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leia" lastname="Fuhrer" birthdate="2012-08-03" gender="F" nation="SUI" license="7175" swrid="5411046" athleteid="12696">
              <RESULTS>
                <RESULT eventid="1068" points="130" swimtime="00:01:47.61" resultid="12697" heatid="14518" lane="3" entrytime="00:01:54.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.77" />
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                    <SPLIT distance="75" swimtime="00:01:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="153" swimtime="00:01:42.52" resultid="12698" heatid="14548" lane="3" entrytime="00:01:40.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.47" />
                    <SPLIT distance="50" swimtime="00:00:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="137" swimtime="00:02:00.74" resultid="12699" heatid="14600" lane="2" entrytime="00:02:02.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.47" />
                    <SPLIT distance="50" swimtime="00:00:58.73" />
                    <SPLIT distance="75" swimtime="00:01:30.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="135" swimtime="00:01:37.78" resultid="12700" heatid="14651" lane="4" entrytime="00:01:35.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.26" />
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="75" swimtime="00:01:11.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yara Jacqueline" lastname="Gfeller" birthdate="2010-01-12" gender="F" nation="SUI" license="7221" swrid="4889115" athleteid="12701">
              <RESULTS>
                <RESULT eventid="1068" points="311" swimtime="00:01:20.54" resultid="12702" heatid="14522" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.98" />
                    <SPLIT distance="50" swimtime="00:00:38.77" />
                    <SPLIT distance="75" swimtime="00:00:59.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="385" swimtime="00:01:15.45" resultid="12703" heatid="14554" lane="2" entrytime="00:01:17.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.59" />
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                    <SPLIT distance="75" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="274" swimtime="00:01:35.95" resultid="12704" heatid="14608" lane="4" entrytime="00:01:38.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.21" />
                    <SPLIT distance="50" swimtime="00:00:45.54" />
                    <SPLIT distance="75" swimtime="00:01:11.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="326" swimtime="00:01:12.99" resultid="12705" heatid="14660" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.70" />
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="75" swimtime="00:00:54.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mara Sophie" lastname="Wiche" birthdate="2011-09-24" gender="F" nation="SUI" license="42335" swrid="5564719" athleteid="12799">
              <RESULTS>
                <RESULT eventid="1078" points="153" swimtime="00:01:42.45" resultid="12800" heatid="14543" lane="4" entrytime="00:01:51.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.97" />
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                    <SPLIT distance="75" swimtime="00:01:18.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="175" swimtime="00:01:51.32" resultid="12801" heatid="14604" lane="2" entrytime="00:01:48.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.25" />
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                    <SPLIT distance="75" swimtime="00:01:21.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="140" swimtime="00:01:36.56" resultid="12802" heatid="14649" lane="3" entrytime="00:01:39.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.68" />
                    <SPLIT distance="50" swimtime="00:00:45.27" />
                    <SPLIT distance="75" swimtime="00:01:12.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konstantinos" lastname="Nath" birthdate="2010-12-28" gender="M" nation="IND" license="42541" swrid="5559275" athleteid="12763">
              <RESULTS>
                <RESULT eventid="1081" points="110" swimtime="00:01:40.79" resultid="12764" heatid="14567" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="97" swimtime="00:02:00.29" resultid="12765" heatid="14621" lane="1" entrytime="00:02:01.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.46" />
                    <SPLIT distance="50" swimtime="00:00:56.38" />
                    <SPLIT distance="75" swimtime="00:01:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="119" swimtime="00:01:31.26" resultid="12766" heatid="14672" lane="3" entrytime="00:01:36.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.01" />
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janis" lastname="Schaller" birthdate="2014-02-07" gender="M" nation="SUI" license="42337" athleteid="12776">
              <RESULTS>
                <RESULT eventid="1066" points="30" swimtime="00:01:09.44" resultid="12777" heatid="14516" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="58" swimtime="00:00:57.11" resultid="12778" heatid="14535" lane="2" entrytime="00:01:01.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="75" swimtime="00:00:47.65" resultid="12779" heatid="14640" lane="4" entrytime="00:00:49.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Léa" lastname="Brechbühler" birthdate="2012-09-15" gender="F" nation="SUI" license="37548" swrid="5484579" athleteid="12688">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende 1) (Zeit: 10:00)" eventid="1078" status="DSQ" swimtime="00:01:49.17" resultid="12689" heatid="14540" lane="2" entrytime="00:02:03.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.94" />
                    <SPLIT distance="50" swimtime="00:00:52.53" />
                    <SPLIT distance="75" swimtime="00:01:19.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="114" swimtime="00:02:08.54" resultid="12690" heatid="14599" lane="3" entrytime="00:02:07.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.76" />
                    <SPLIT distance="50" swimtime="00:01:00.54" />
                    <SPLIT distance="75" swimtime="00:01:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="148" swimtime="00:01:34.96" resultid="12691" heatid="14647" lane="3" entrytime="00:01:44.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.64" />
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="75" swimtime="00:01:10.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandros" lastname="Kokkalis" birthdate="2010-04-22" gender="M" nation="SUI" license="7123" swrid="5244624" athleteid="12725">
              <RESULTS>
                <RESULT eventid="1071" points="86" swimtime="00:01:48.24" resultid="12726" heatid="14525" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.24" />
                    <SPLIT distance="50" swimtime="00:00:47.77" />
                    <SPLIT distance="75" swimtime="00:01:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="172" swimtime="00:01:26.75" resultid="12727" heatid="14571" lane="2" entrytime="00:01:30.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.11" />
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="186" swimtime="00:01:36.79" resultid="12728" heatid="14628" lane="2" entrytime="00:01:36.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.72" />
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                    <SPLIT distance="75" swimtime="00:01:11.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="211" swimtime="00:01:15.41" resultid="12729" heatid="14680" lane="1" entrytime="00:01:15.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.19" />
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                    <SPLIT distance="75" swimtime="00:00:56.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elin" lastname="Schwab" birthdate="2011-01-24" gender="F" nation="SUI" license="7148" swrid="5335433" athleteid="12785">
              <RESULTS>
                <RESULT eventid="1068" points="161" swimtime="00:01:40.32" resultid="12786" heatid="14520" lane="4" entrytime="00:01:42.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.41" />
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                    <SPLIT distance="75" swimtime="00:01:12.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="204" swimtime="00:01:33.15" resultid="12787" heatid="14551" lane="4" entrytime="00:01:35.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:10.34" />
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="183" swimtime="00:01:49.65" resultid="12788" heatid="14603" lane="3" entrytime="00:01:50.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.53" />
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                    <SPLIT distance="75" swimtime="00:01:20.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="230" swimtime="00:01:22.00" resultid="12789" heatid="14655" lane="2" entrytime="00:01:24.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.50" />
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="75" swimtime="00:01:01.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nikos" lastname="Kokkalis" birthdate="2012-04-27" gender="M" nation="SUI" license="7198" swrid="5335428" athleteid="12730">
              <RESULTS>
                <RESULT eventid="1081" points="107" swimtime="00:01:41.53" resultid="12731" heatid="14567" lane="3" entrytime="00:01:45.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.67" />
                    <SPLIT distance="50" swimtime="00:00:50.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="119" swimtime="00:01:52.25" resultid="12732" heatid="14620" lane="3" entrytime="00:02:04.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.55" />
                    <SPLIT distance="50" swimtime="00:00:53.73" />
                    <SPLIT distance="75" swimtime="00:01:23.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="124" swimtime="00:01:29.90" resultid="12733" heatid="14675" lane="3" entrytime="00:01:31.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.00" />
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="75" swimtime="00:01:06.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luc" lastname="Willen" birthdate="2010-12-12" gender="M" nation="SUI" license="7187" swrid="5387430" athleteid="12807">
              <RESULTS>
                <RESULT eventid="1071" points="156" swimtime="00:01:28.68" resultid="12808" heatid="14526" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.80" />
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                    <SPLIT distance="75" swimtime="00:01:01.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="212" swimtime="00:01:20.94" resultid="12809" heatid="14573" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="75" swimtime="00:01:01.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="208" swimtime="00:01:33.32" resultid="12810" heatid="14629" lane="1" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.27" />
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                    <SPLIT distance="75" swimtime="00:01:08.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="246" swimtime="00:01:11.65" resultid="12811" heatid="14681" lane="3" entrytime="00:01:09.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.90" />
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="75" swimtime="00:00:53.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryan" lastname="Rybarczyk" birthdate="2014-03-06" gender="M" nation="SUI" license="40492" swrid="5509064" athleteid="12772">
              <RESULTS>
                <RESULT eventid="1076" points="74" swimtime="00:00:52.75" resultid="12773" heatid="14537" lane="4" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="78" swimtime="00:00:59.07" resultid="12774" heatid="14592" lane="2" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="65" swimtime="00:00:50.11" resultid="12775" heatid="14640" lane="1" entrytime="00:00:49.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lisa" lastname="Leupi" birthdate="2010-08-31" gender="F" nation="SUI" license="7182" swrid="5243021" athleteid="12742">
              <RESULTS>
                <RESULT eventid="1068" points="276" swimtime="00:01:23.84" resultid="12743" heatid="14522" lane="2" entrytime="00:01:21.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.46" />
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="75" swimtime="00:01:01.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="339" swimtime="00:01:18.69" resultid="12744" heatid="14554" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.30" />
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                    <SPLIT distance="75" swimtime="00:00:58.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="275" swimtime="00:01:35.89" resultid="12745" heatid="14609" lane="3" entrytime="00:01:34.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.09" />
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="75" swimtime="00:01:11.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="344" swimtime="00:01:11.68" resultid="12746" heatid="14660" lane="2" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.53" />
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauryn" lastname="Ghiggia" birthdate="2011-10-10" gender="F" nation="SUI" license="7172" swrid="5411040" athleteid="12706">
              <RESULTS>
                <RESULT eventid="1092" points="285" swimtime="00:01:34.66" resultid="12707" heatid="14608" lane="1" entrytime="00:01:37.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.26" />
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="75" swimtime="00:01:09.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="209" swimtime="00:01:24.56" resultid="12708" heatid="14656" lane="3" entrytime="00:01:23.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.95" />
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="75" swimtime="00:01:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="168" swimtime="00:01:38.89" resultid="12709" heatid="14520" lane="2" entrytime="00:01:37.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.34" />
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="75" swimtime="00:01:12.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="201" swimtime="00:01:33.61" resultid="12710" heatid="14549" lane="4" entrytime="00:01:38.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.02" />
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="75" swimtime="00:01:09.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Silian Lias" lastname="Gschwend" birthdate="2010-06-21" gender="M" nation="SUI" license="7212" swrid="5326500" athleteid="12711">
              <RESULTS>
                <RESULT eventid="1071" points="144" swimtime="00:01:31.02" resultid="12712" heatid="14526" lane="1" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.17" />
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="75" swimtime="00:01:05.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="196" swimtime="00:01:23.17" resultid="12713" heatid="14573" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.42" />
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="75" swimtime="00:01:03.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="258" swimtime="00:01:26.88" resultid="12714" heatid="14629" lane="2" entrytime="00:01:27.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.37" />
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="75" swimtime="00:01:04.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="225" swimtime="00:01:13.84" resultid="12715" heatid="14681" lane="4" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.17" />
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="75" swimtime="00:00:55.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dario" lastname="Meier" birthdate="2011-08-22" gender="M" nation="SUI" license="27425" swrid="5464178" athleteid="12751">
              <RESULTS>
                <RESULT eventid="1081" points="88" swimtime="00:01:48.44" resultid="12752" heatid="14569" lane="3" entrytime="00:01:40.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.63" />
                    <SPLIT distance="50" swimtime="00:00:51.13" />
                    <SPLIT distance="75" swimtime="00:01:20.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="139" swimtime="00:01:46.70" resultid="12753" heatid="14625" lane="2" entrytime="00:01:49.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.47" />
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                    <SPLIT distance="75" swimtime="00:01:17.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="129" swimtime="00:01:28.79" resultid="12754" heatid="14676" lane="2" entrytime="00:01:28.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.12" />
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                    <SPLIT distance="75" swimtime="00:01:05.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmina" lastname="Melotte" birthdate="2011-07-08" gender="F" nation="SUI" license="27780" swrid="5467815" athleteid="12755">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="12756" entrytime="00:01:44.78" entrycourse="SCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="12757" entrytime="00:01:55.51" entrycourse="SCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="12758" entrytime="00:01:31.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lennox" lastname="Sutter" birthdate="2012-08-22" gender="M" nation="SUI" license="7176" swrid="5411052" athleteid="12795">
              <RESULTS>
                <RESULT eventid="1081" points="138" swimtime="00:01:33.49" resultid="12796" heatid="14571" lane="4" entrytime="00:01:33.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.16" />
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="206 - Unterwasserphase: Mehr als ein Delphinbeinschlag (Start) (Zeit: 13:24)" eventid="1095" status="DSQ" swimtime="00:01:44.60" resultid="12797" heatid="14628" lane="4" entrytime="00:01:41.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.99" />
                    <SPLIT distance="50" swimtime="00:00:49.57" />
                    <SPLIT distance="75" swimtime="00:01:18.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="121" swimtime="00:01:30.77" resultid="12798" heatid="14678" lane="4" entrytime="00:01:25.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.80" />
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="75" swimtime="00:01:08.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jonas" lastname="Leupi" birthdate="2012-07-01" gender="M" nation="SUI" license="7186" swrid="5411043" athleteid="12738">
              <RESULTS>
                <RESULT eventid="1081" points="84" swimtime="00:01:50.04" resultid="12739" heatid="14566" lane="3" entrytime="00:01:48.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="90" swimtime="00:02:03.42" resultid="12740" heatid="14617" lane="3" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.06" />
                    <SPLIT distance="50" swimtime="00:01:00.47" />
                    <SPLIT distance="75" swimtime="00:01:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="96" swimtime="00:01:37.89" resultid="12741" heatid="14674" lane="4" entrytime="00:01:34.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                    <SPLIT distance="75" swimtime="00:01:14.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Annik" lastname="Maurer" birthdate="2011-07-14" gender="F" nation="SUI" license="7128" swrid="5353512" athleteid="12747">
              <RESULTS>
                <RESULT eventid="1078" points="205" swimtime="00:01:33.08" resultid="12748" heatid="14550" lane="3" entrytime="00:01:36.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.34" />
                    <SPLIT distance="50" swimtime="00:00:45.44" />
                    <SPLIT distance="75" swimtime="00:01:09.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="171" swimtime="00:01:52.30" resultid="12749" heatid="14603" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.79" />
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                    <SPLIT distance="75" swimtime="00:01:23.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="217" swimtime="00:01:23.59" resultid="12750" heatid="14654" lane="2" entrytime="00:01:25.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.46" />
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                    <SPLIT distance="75" swimtime="00:01:02.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yul" lastname="Rüfenacht" birthdate="2010-01-21" gender="M" nation="SUI" license="7222" swrid="5243039" athleteid="12767">
              <RESULTS>
                <RESULT eventid="1071" points="86" swimtime="00:01:48.19" resultid="12768" heatid="14525" lane="4" entrytime="00:01:51.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="150" swimtime="00:01:30.95" resultid="12769" heatid="14572" lane="3" entrytime="00:01:28.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.60" />
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                    <SPLIT distance="75" swimtime="00:01:08.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="139" swimtime="00:01:46.71" resultid="12770" heatid="14627" lane="1" entrytime="00:01:43.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.16" />
                    <SPLIT distance="50" swimtime="00:00:50.04" />
                    <SPLIT distance="75" swimtime="00:01:19.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="150" swimtime="00:01:24.52" resultid="12771" heatid="14679" lane="1" entrytime="00:01:19.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.59" />
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="75" swimtime="00:01:02.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aurelia" lastname="Scheurer" birthdate="2011-01-16" gender="F" nation="SUI" license="7130" swrid="5335438" athleteid="12780">
              <RESULTS>
                <RESULT eventid="1068" points="257" swimtime="00:01:25.81" resultid="12781" heatid="14521" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.74" />
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="75" swimtime="00:01:02.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="303" swimtime="00:01:21.66" resultid="12782" heatid="14554" lane="1" entrytime="00:01:18.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.12" />
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="75" swimtime="00:01:01.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="348" swimtime="00:01:28.59" resultid="12783" heatid="14610" lane="3" entrytime="00:01:28.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.73" />
                    <SPLIT distance="50" swimtime="00:00:41.71" />
                    <SPLIT distance="75" swimtime="00:01:05.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="372" swimtime="00:01:09.83" resultid="12784" heatid="14660" lane="1" entrytime="00:01:12.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.09" />
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="75" swimtime="00:00:52.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noemi" lastname="Wichtermann" birthdate="2011-10-17" gender="F" nation="SUI" license="35796" swrid="5484577" athleteid="12803">
              <RESULTS>
                <RESULT eventid="1078" points="117" swimtime="00:01:51.99" resultid="12804" heatid="14542" lane="4" entrytime="00:01:58.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.10" />
                    <SPLIT distance="50" swimtime="00:00:56.44" />
                    <SPLIT distance="75" swimtime="00:01:25.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="142" swimtime="00:01:59.40" resultid="12805" heatid="14598" lane="2" entrytime="00:02:09.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.00" />
                    <SPLIT distance="50" swimtime="00:00:56.18" />
                    <SPLIT distance="75" swimtime="00:01:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="105" swimtime="00:01:46.22" resultid="12806" heatid="14645" lane="4" entrytime="00:02:03.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.15" />
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                    <SPLIT distance="75" swimtime="00:01:20.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yousra" lastname="Berrichi" birthdate="2012-05-15" gender="F" nation="FRA" license="32121" swrid="5464133" athleteid="12683">
              <RESULTS>
                <RESULT eventid="1068" points="122" swimtime="00:01:49.86" resultid="12684" heatid="14519" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.46" />
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                    <SPLIT distance="75" swimtime="00:01:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="232" swimtime="00:01:29.21" resultid="12685" heatid="14552" lane="3" entrytime="00:01:32.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="191" swimtime="00:01:48.27" resultid="12686" heatid="14605" lane="1" entrytime="00:01:45.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.01" />
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                    <SPLIT distance="75" swimtime="00:01:19.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="224" swimtime="00:01:22.73" resultid="12687" heatid="14655" lane="1" entrytime="00:01:25.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.30" />
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="75" swimtime="00:01:02.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erik" lastname="Hirsbrunner" birthdate="2011-07-09" gender="M" nation="SUI" license="32138" swrid="5464168" athleteid="12716">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende 1) (Zeit: 10:47)" eventid="1081" status="DSQ" swimtime="00:01:37.03" resultid="12717" heatid="14569" lane="2" entrytime="00:01:38.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.20" />
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="75" swimtime="00:01:12.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="92" swimtime="00:02:02.57" resultid="12718" heatid="14620" lane="2" entrytime="00:02:03.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.36" />
                    <SPLIT distance="50" swimtime="00:00:57.67" />
                    <SPLIT distance="75" swimtime="00:01:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="153" swimtime="00:01:23.85" resultid="12719" heatid="14678" lane="1" entrytime="00:01:24.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.35" />
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="75" swimtime="00:01:01.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Saga" lastname="Hirsbrunner" birthdate="2013-08-26" gender="F" nation="SUI" license="37458" swrid="5484581" athleteid="12720">
              <RESULTS>
                <RESULT eventid="1064" points="86" swimtime="00:00:55.08" resultid="12721" heatid="14514" lane="2" entrytime="00:00:55.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="160" swimtime="00:00:47.12" resultid="12722" heatid="14533" lane="4" entrytime="00:00:48.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="145" swimtime="00:00:54.25" resultid="12723" heatid="14588" lane="2" entrytime="00:00:59.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="171" swimtime="00:00:41.29" resultid="12724" heatid="14637" lane="4" entrytime="00:00:41.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="231" swimtime="00:02:13.25" resultid="12817" heatid="14818" lane="2" entrytime="00:02:13.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="75" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="125" swimtime="00:01:22.17" />
                    <SPLIT distance="150" swimtime="00:01:39.44" />
                    <SPLIT distance="175" swimtime="00:01:55.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12711" number="1" />
                    <RELAYPOSITION athleteid="12807" number="2" />
                    <RELAYPOSITION athleteid="12790" number="3" />
                    <RELAYPOSITION athleteid="12725" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer 2) (Zeit: 11:34)" eventid="1086" status="DSQ" swimtime="00:02:30.78" resultid="12818" heatid="14583" lane="2" entrytime="00:02:26.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="75" swimtime="00:00:53.67" />
                    <SPLIT distance="100" swimtime="00:01:14.75" />
                    <SPLIT distance="125" swimtime="00:01:31.63" />
                    <SPLIT distance="150" swimtime="00:01:50.54" />
                    <SPLIT distance="175" swimtime="00:02:10.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12767" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="12763" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="12716" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="12734" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="3">
              <RESULTS>
                <RESULT eventid="1086" points="127" swimtime="00:02:42.38" resultid="12819" heatid="14583" lane="4" entrytime="00:02:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.46" />
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="75" swimtime="00:00:59.78" />
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="125" swimtime="00:01:39.26" />
                    <SPLIT distance="150" swimtime="00:02:01.20" />
                    <SPLIT distance="175" swimtime="00:02:20.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12759" number="1" />
                    <RELAYPOSITION athleteid="12795" number="2" />
                    <RELAYPOSITION athleteid="12730" number="3" />
                    <RELAYPOSITION athleteid="12738" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="4">
              <RESULTS>
                <RESULT eventid="1086" points="94" status="EXH" swimtime="00:02:59.47" resultid="12820" heatid="14581" lane="1" entrytime="00:03:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.50" />
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="75" swimtime="00:01:03.02" />
                    <SPLIT distance="100" swimtime="00:01:29.95" />
                    <SPLIT distance="125" swimtime="00:01:51.65" />
                    <SPLIT distance="150" swimtime="00:02:15.23" />
                    <SPLIT distance="175" swimtime="00:02:34.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12751" number="1" />
                    <RELAYPOSITION athleteid="12772" number="2" />
                    <RELAYPOSITION athleteid="12776" number="3" />
                    <RELAYPOSITION athleteid="12688" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="378" swimtime="00:02:07.90" resultid="12821" heatid="14817" lane="3" entrytime="00:02:11.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="75" swimtime="00:00:47.74" />
                    <SPLIT distance="100" swimtime="00:01:04.53" />
                    <SPLIT distance="125" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:01:36.88" />
                    <SPLIT distance="175" swimtime="00:01:51.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12812" number="1" />
                    <RELAYPOSITION athleteid="12701" number="2" />
                    <RELAYPOSITION athleteid="12742" number="3" />
                    <RELAYPOSITION athleteid="12780" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1084" points="235" swimtime="00:02:29.81" resultid="12822" heatid="14817" lane="4" entrytime="00:02:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.83" />
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="75" swimtime="00:00:53.26" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="125" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                    <SPLIT distance="175" swimtime="00:02:07.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12683" number="1" />
                    <RELAYPOSITION athleteid="12706" number="2" />
                    <RELAYPOSITION athleteid="12785" number="3" />
                    <RELAYPOSITION athleteid="12696" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1084" points="158" swimtime="00:02:50.76" resultid="12823" heatid="14578" lane="2" entrytime="00:02:44.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="75" swimtime="00:00:59.02" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="125" swimtime="00:01:43.58" />
                    <SPLIT distance="150" swimtime="00:02:05.46" />
                    <SPLIT distance="175" swimtime="00:02:27.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12747" number="1" />
                    <RELAYPOSITION athleteid="12720" number="2" />
                    <RELAYPOSITION athleteid="12799" number="3" />
                    <RELAYPOSITION athleteid="12803" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="TAGI" nation="SUI" region="RZO" clubid="13243" swrid="65626" name="Schwimmclub Tägi Wettingen">
          <ATHLETES>
            <ATHLETE firstname="Stella" lastname="Schneider" birthdate="2011-01-31" gender="F" nation="SUI" swrid="5489043" athleteid="13318">
              <RESULTS>
                <RESULT eventid="1092" points="240" swimtime="00:01:40.26" resultid="13319" heatid="14602" lane="2" entrytime="00:01:52.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.80" />
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="75" swimtime="00:01:10.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="223" swimtime="00:01:22.80" resultid="13320" heatid="14651" lane="3" entrytime="00:01:34.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                    <SPLIT distance="75" swimtime="00:01:00.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucia" lastname="Bermudez - Casal" birthdate="2010-10-04" gender="F" nation="ESP" swrid="5419928" athleteid="13244">
              <RESULTS>
                <RESULT eventid="1078" points="182" swimtime="00:01:36.76" resultid="13245" heatid="14544" lane="1" entrytime="00:01:48.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.48" />
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                    <SPLIT distance="75" swimtime="00:01:11.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="212" swimtime="00:01:24.16" resultid="13246" heatid="14656" lane="2" entrytime="00:01:23.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luna" lastname="Buchser" birthdate="2011-07-17" gender="F" nation="SUI" athleteid="13265">
              <RESULTS>
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="13266" entrytime="00:01:42.07" entrycourse="SCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13267" entrytime="00:01:58.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rebecca" lastname="Neuberth" birthdate="2009-01-31" gender="F" nation="SUI" swrid="5489040" athleteid="13304">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="13305" entrytime="00:01:33.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Seraina" lastname="Kaup" birthdate="2009-06-23" gender="F" nation="SUI" license="119442" swrid="5326620" athleteid="13286">
              <RESULTS>
                <RESULT eventid="1114" points="249" swimtime="00:01:27.16" resultid="13287" heatid="14707" lane="4" entrytime="00:01:28.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="75" swimtime="00:01:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="262" swimtime="00:01:18.48" resultid="13288" heatid="14768" lane="1" entrytime="00:01:19.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.86" />
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                    <SPLIT distance="75" swimtime="00:00:58.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tilia" lastname="Hil" birthdate="2006-07-25" gender="F" nation="AUT" license="103951" swrid="5053816" athleteid="13280">
              <RESULTS>
                <RESULT eventid="1124" points="278" swimtime="00:01:35.50" resultid="13281" heatid="14742" lane="2" entrytime="00:01:35.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.75" />
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                    <SPLIT distance="75" swimtime="00:01:10.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="295" swimtime="00:01:15.45" resultid="13282" heatid="14769" lane="2" entrytime="00:01:15.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.41" />
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="75" swimtime="00:00:56.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolin" lastname="Hil" birthdate="2011-11-17" gender="F" nation="SUI" swrid="5298337" athleteid="13277">
              <RESULTS>
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13278" entrytime="00:02:05.00" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="13279" entrytime="00:01:44.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Rutz" birthdate="2010-09-21" gender="F" nation="SUI" athleteid="13312">
              <RESULTS>
                <RESULT eventid="1102" points="143" swimtime="00:01:35.97" resultid="13313" heatid="14648" lane="3" entrytime="00:01:41.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="136" swimtime="00:01:46.60" resultid="13314" heatid="14543" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.85" />
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="75" swimtime="00:01:18.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuel" lastname="Simeoni" birthdate="2005-08-27" gender="M" nation="SUI" license="104778" swrid="5068074" athleteid="13321">
              <RESULTS>
                <RESULT comment="999 - , eigene Bahn verlassen" eventid="1117" status="DSQ" swimtime="00:01:15.60" resultid="13322" heatid="14726" lane="2" entrytime="00:01:09.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.77" />
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="441" swimtime="00:00:59.02" resultid="13323" heatid="14793" lane="1" entrytime="00:00:59.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Bozinov" birthdate="2010-03-26" gender="M" nation="MKD" license="119042" swrid="5314584" athleteid="13259">
              <RESULTS>
                <RESULT eventid="1081" points="170" swimtime="00:01:27.10" resultid="13260" heatid="14571" lane="1" entrytime="00:01:33.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.87" />
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="229" swimtime="00:01:13.37" resultid="13261" heatid="14680" lane="3" entrytime="00:01:15.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.06" />
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="75" swimtime="00:00:54.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elin" lastname="Buchser" birthdate="2012-09-04" gender="F" nation="SUI" athleteid="13262">
              <RESULTS>
                <RESULT eventid="1102" points="96" swimtime="00:01:49.71" resultid="13263" heatid="14644" lane="2" entrytime="00:02:08.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:24.58" />
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="144" swimtime="00:01:58.93" resultid="13264" heatid="14596" lane="1" entrytime="00:02:22.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.34" />
                    <SPLIT distance="50" swimtime="00:00:56.46" />
                    <SPLIT distance="75" swimtime="00:01:29.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alicia" lastname="Meta" birthdate="2010-11-11" gender="F" nation="SUI" swrid="5489038" athleteid="13301">
              <RESULTS>
                <RESULT eventid="1078" points="134" swimtime="00:01:47.11" resultid="13302" heatid="14545" lane="2" entrytime="00:01:45.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.99" />
                    <SPLIT distance="50" swimtime="00:00:51.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="213" swimtime="00:01:24.02" resultid="13303" heatid="14655" lane="4" entrytime="00:01:25.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.76" />
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="75" swimtime="00:01:02.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daphne" lastname="Passmore" birthdate="2012-01-02" gender="F" nation="SUI" athleteid="13306">
              <RESULTS>
                <RESULT eventid="1102" points="115" swimtime="00:01:43.18" resultid="13307" heatid="14649" lane="4" entrytime="00:01:39.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="139" swimtime="00:01:45.77" resultid="13308" heatid="14543" lane="3" entrytime="00:01:51.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.37" />
                    <SPLIT distance="50" swimtime="00:00:48.61" />
                    <SPLIT distance="75" swimtime="00:01:17.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leena" lastname="Kosonen" birthdate="2012-06-19" gender="F" nation="SUI" athleteid="13292">
              <RESULTS>
                <RESULT comment="302 - Wand nicht berührt (Wende ...) (Zeit: 9:56)" eventid="1078" status="DSQ" swimtime="00:02:12.21" resultid="13293" heatid="14539" lane="4" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.05" />
                    <SPLIT distance="75" swimtime="00:01:40.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="82" swimtime="00:01:55.50" resultid="13294" heatid="14645" lane="1" entrytime="00:02:00.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.40" />
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                    <SPLIT distance="75" swimtime="00:01:26.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jules" lastname="Hübscher" birthdate="2012-09-23" gender="M" nation="SUI" swrid="5301986" athleteid="13283">
              <RESULTS>
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="13284" entrytime="00:02:00.00" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="13285" entrytime="00:01:38.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ella" lastname="Bouvard" birthdate="2009-12-11" gender="F" nation="SUI" swrid="5489033" athleteid="13253">
              <RESULTS>
                <RESULT eventid="1108" points="320" swimtime="00:01:19.83" resultid="13254" heatid="14686" lane="2" entrytime="00:01:28.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.56" />
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="75" swimtime="00:00:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="352" swimtime="00:01:11.13" resultid="13255" heatid="14770" lane="3" entrytime="00:01:14.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.97" />
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="75" swimtime="00:00:52.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Levi" lastname="Bouvard" birthdate="2011-06-28" gender="M" nation="SUI" swrid="5489034" athleteid="13256">
              <RESULTS>
                <RESULT eventid="1095" points="150" swimtime="00:01:44.09" resultid="13257" heatid="14626" lane="3" entrytime="00:01:47.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.84" />
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                    <SPLIT distance="75" swimtime="00:01:17.84" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 14:47)" eventid="1105" status="DSQ" swimtime="00:01:23.48" resultid="13258" heatid="14675" lane="1" entrytime="00:01:32.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.67" />
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="75" swimtime="00:01:03.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Janick" lastname="Zimmerli" birthdate="2001-12-03" gender="M" nation="SUI" license="29706" swrid="4781061" athleteid="13330">
              <RESULTS>
                <RESULT eventid="1111" points="546" swimtime="00:00:58.45" resultid="13331" heatid="14701" lane="4" entrytime="00:00:59.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.48" />
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                    <SPLIT distance="75" swimtime="00:00:42.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="525" swimtime="00:00:55.70" resultid="13332" heatid="14795" lane="3" entrytime="00:00:56.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:26.82" />
                    <SPLIT distance="75" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="460" swimtime="00:00:28.77" resultid="14859" heatid="14843" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="My-An" lastname="Lauber" birthdate="2010-02-01" gender="F" nation="SUI" swrid="5489037" athleteid="13295">
              <RESULTS>
                <RESULT eventid="1092" points="262" swimtime="00:01:37.43" resultid="13296" heatid="14609" lane="2" entrytime="00:01:32.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.20" />
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="75" swimtime="00:01:10.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="229" swimtime="00:01:22.05" resultid="13297" heatid="14655" lane="3" entrytime="00:01:24.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.29" />
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="75" swimtime="00:00:59.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlon" lastname="Umbricht" birthdate="2013-01-23" gender="M" nation="SUI" athleteid="13327">
              <RESULTS>
                <RESULT eventid="1100" points="111" swimtime="00:00:41.86" resultid="13328" heatid="14641" lane="4" entrytime="00:00:45.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="85" swimtime="00:00:57.29" resultid="13329" heatid="14593" lane="3" entrytime="00:01:02.88">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leano" lastname="Schmid" birthdate="2010-10-09" gender="M" nation="SUI" swrid="5489042" athleteid="13315">
              <RESULTS>
                <RESULT eventid="1095" points="155" swimtime="00:01:42.81" resultid="13316" heatid="14627" lane="3" entrytime="00:01:43.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.65" />
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                    <SPLIT distance="75" swimtime="00:01:14.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="129" swimtime="00:01:28.91" resultid="13317" heatid="14676" lane="3" entrytime="00:01:29.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.33" />
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="75" swimtime="00:01:06.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Del Toro" birthdate="2008-05-15" gender="F" nation="SUI" license="119047" swrid="5314586" athleteid="13268">
              <RESULTS>
                <RESULT eventid="1114" points="183" swimtime="00:01:36.56" resultid="13269" heatid="14704" lane="1" entrytime="00:01:45.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="277" swimtime="00:01:17.04" resultid="13270" heatid="14768" lane="4" entrytime="00:01:20.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="75" swimtime="00:00:57.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Gysel" birthdate="2008-02-25" gender="F" nation="SUI" license="109957" swrid="5178021" athleteid="13272">
              <RESULTS>
                <RESULT eventid="1124" points="300" swimtime="00:01:33.15" resultid="13273" heatid="14744" lane="4" entrytime="00:01:32.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.09" />
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="75" swimtime="00:01:08.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelie" lastname="Hil" birthdate="2009-11-09" gender="F" nation="SUI" license="119046" swrid="5314587" athleteid="13274">
              <RESULTS>
                <RESULT eventid="1124" points="273" swimtime="00:01:36.08" resultid="13275" heatid="14742" lane="3" entrytime="00:01:35.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.88" />
                    <SPLIT distance="50" swimtime="00:00:45.51" />
                    <SPLIT distance="75" swimtime="00:01:10.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="279" swimtime="00:01:16.89" resultid="13276" heatid="14768" lane="3" entrytime="00:01:19.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="75" swimtime="00:00:57.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristina" lastname="Eichenberger" birthdate="2008-05-12" gender="F" nation="SUI" license="109958" swrid="5083241" athleteid="13271" />
            <ATHLETE firstname="My-Son" lastname="Lauber" birthdate="2012-06-11" gender="M" nation="SUI" athleteid="13298">
              <RESULTS>
                <RESULT eventid="1105" points="102" swimtime="00:01:36.15" resultid="13299" heatid="14672" lane="2" entrytime="00:01:36.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.32" />
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="75" swimtime="00:01:10.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="93" swimtime="00:02:01.99" resultid="13300" heatid="14625" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.48" />
                    <SPLIT distance="50" swimtime="00:00:57.31" />
                    <SPLIT distance="75" swimtime="00:01:30.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Bolliger" birthdate="2007-06-24" gender="M" nation="SUI" license="121518" swrid="5353381" athleteid="13250">
              <RESULTS>
                <RESULT eventid="1117" points="215" swimtime="00:01:20.66" resultid="13251" heatid="14721" lane="2" entrytime="00:01:25.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.99" />
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="75" swimtime="00:00:59.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="330" swimtime="00:01:05.02" resultid="13252" heatid="14790" lane="1" entrytime="00:01:04.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.90" />
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="75" swimtime="00:00:48.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Stommel Minamisawa" birthdate="2013-10-24" gender="M" nation="GER" athleteid="13324">
              <RESULTS>
                <RESULT eventid="1090" points="70" swimtime="00:01:01.24" resultid="13325" heatid="14593" lane="1" entrytime="00:01:03.38">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="81" swimtime="00:00:46.55" resultid="13326" heatid="14639" lane="3" entrytime="00:00:53.27" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nada" lastname="Klaric" birthdate="2007-09-08" gender="F" nation="SUI" athleteid="13289">
              <RESULTS>
                <RESULT eventid="1108" points="312" swimtime="00:01:20.47" resultid="13290" heatid="14686" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="75" swimtime="00:00:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="389" swimtime="00:01:08.83" resultid="13291" heatid="14773" lane="4" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.05" />
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                    <SPLIT distance="75" swimtime="00:00:50.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrei" lastname="Bertea" birthdate="2006-10-27" gender="M" nation="SUI" license="36781" swrid="5299844" athleteid="13247">
              <RESULTS>
                <RESULT eventid="1127" points="316" swimtime="00:01:21.18" resultid="13248" heatid="14759" lane="3" entrytime="00:01:23.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.40" />
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                    <SPLIT distance="75" swimtime="00:00:59.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="304" swimtime="00:01:06.82" resultid="13249" heatid="14789" lane="1" entrytime="00:01:06.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.44" />
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="75" swimtime="00:00:50.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Robertson" birthdate="2011-10-16" gender="F" nation="AUS" swrid="5489041" athleteid="13309">
              <RESULTS>
                <RESULT comment="999 - , 209 Zehen beim Start nicht an der Wand" eventid="1078" status="DSQ" swimtime="00:01:47.04" resultid="13310" heatid="14542" lane="1" entrytime="00:01:56.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.25" />
                    <SPLIT distance="50" swimtime="00:00:51.21" />
                    <SPLIT distance="75" swimtime="00:01:20.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="193" swimtime="00:01:26.85" resultid="13311" heatid="14652" lane="3" entrytime="00:01:30.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.93" />
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="75" swimtime="00:01:04.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="146" swimtime="00:02:35.22" resultid="13333" heatid="14582" lane="2" entrytime="00:02:43.34">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.74" />
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="75" swimtime="00:00:52.52" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="125" swimtime="00:01:35.78" />
                    <SPLIT distance="150" swimtime="00:01:58.61" />
                    <SPLIT distance="175" swimtime="00:02:16.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13259" number="1" />
                    <RELAYPOSITION athleteid="13315" number="2" />
                    <RELAYPOSITION athleteid="13327" number="3" />
                    <RELAYPOSITION athleteid="13256" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="384" swimtime="00:02:04.32" resultid="13334" heatid="14736" lane="4" entrytime="00:02:05.43">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.72" />
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="75" swimtime="00:00:52.18" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="125" swimtime="00:01:24.00" />
                    <SPLIT distance="150" swimtime="00:01:38.27" />
                    <SPLIT distance="175" swimtime="00:01:50.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13250" number="1" />
                    <RELAYPOSITION athleteid="13247" number="2" />
                    <RELAYPOSITION athleteid="13330" number="3" />
                    <RELAYPOSITION athleteid="13321" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="243" swimtime="00:02:28.15" resultid="13335" heatid="14579" lane="1" entrytime="00:02:39.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.85" />
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="75" swimtime="00:00:54.57" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="125" swimtime="00:01:32.56" />
                    <SPLIT distance="150" swimtime="00:01:51.73" />
                    <SPLIT distance="175" swimtime="00:02:09.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13244" number="1" />
                    <RELAYPOSITION athleteid="13301" number="2" />
                    <RELAYPOSITION athleteid="13318" number="3" />
                    <RELAYPOSITION athleteid="13295" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="303" swimtime="00:02:32.29" resultid="13336" heatid="14731" lane="1" entrytime="00:02:38.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="75" swimtime="00:00:58.61" />
                    <SPLIT distance="100" swimtime="00:01:21.88" />
                    <SPLIT distance="125" swimtime="00:01:38.00" />
                    <SPLIT distance="150" swimtime="00:01:57.23" />
                    <SPLIT distance="175" swimtime="00:02:14.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13253" number="1" />
                    <RELAYPOSITION athleteid="13280" number="2" />
                    <RELAYPOSITION athleteid="13289" number="3" />
                    <RELAYPOSITION athleteid="13268" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1084" points="125" swimtime="00:03:04.82" resultid="13337" heatid="14577" lane="3" entrytime="00:03:04.19">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.28" />
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                    <SPLIT distance="75" swimtime="00:01:14.19" />
                    <SPLIT distance="100" swimtime="00:01:41.83" />
                    <SPLIT distance="125" swimtime="00:02:01.64" />
                    <SPLIT distance="150" swimtime="00:02:23.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13262" number="1" />
                    <RELAYPOSITION athleteid="13292" number="2" />
                    <RELAYPOSITION athleteid="13312" number="3" />
                    <RELAYPOSITION athleteid="13309" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1120" status="WDR" swimtime="00:00:00.00" resultid="13338" entrytime="00:02:55.40">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13286" number="1" />
                    <RELAYPOSITION athleteid="13280" number="2" />
                    <RELAYPOSITION athleteid="13274" number="3" />
                    <RELAYPOSITION athleteid="13268" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BAAR" nation="SUI" region="RZO" clubid="13981" swrid="65640" name="Schwimmverein Baar" shortname="SV Baar">
          <ATHLETES>
            <ATHLETE firstname="Leo" lastname="Verschooten" birthdate="2006-03-26" gender="M" nation="BEL" license="119231" swrid="5314511" athleteid="13985" level="INT/NAT">
              <RESULTS>
                <RESULT eventid="1127" points="479" swimtime="00:01:10.71" resultid="13986" heatid="14762" lane="2" entrytime="00:01:07.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.81" />
                    <SPLIT distance="50" swimtime="00:00:32.80" />
                    <SPLIT distance="75" swimtime="00:00:51.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="600" swimtime="00:00:53.28" resultid="13987" heatid="14797" lane="2" entrytime="00:00:51.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.89" />
                    <SPLIT distance="50" swimtime="00:00:24.99" />
                    <SPLIT distance="75" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="545" swimtime="00:00:27.20" resultid="14858" heatid="14843" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6683" points="487" swimtime="00:00:32.08" resultid="14868" heatid="14804" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6639" points="603" swimtime="00:00:25.74" resultid="14873" heatid="14806" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6679" points="624" swimtime="00:00:23.58" resultid="14878" heatid="14808" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mia-Lena" lastname="Sigrist" birthdate="2007-01-13" gender="F" nation="SUI" license="111710" swrid="4821638" athleteid="13982" level="KSK/RZO">
              <RESULTS>
                <RESULT eventid="1124" points="504" swimtime="00:01:18.33" resultid="13983" heatid="14750" lane="3" entrytime="00:01:14.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.23" />
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="75" swimtime="00:00:57.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="493" swimtime="00:01:03.58" resultid="13984" heatid="14780" lane="1" entrytime="00:01:01.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.34" />
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="75" swimtime="00:00:46.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WSCK" nation="SUI" region="RZO" clubid="12597" swrid="65644" name="Wassersport-Club Kloten">
          <ATHLETES>
            <ATHLETE firstname="Massimo" lastname="Rossi" birthdate="2007-01-27" gender="M" nation="SUI" license="8025" swrid="5150421" athleteid="12645">
              <RESULTS>
                <RESULT eventid="1117" points="332" swimtime="00:01:09.76" resultid="12646" heatid="14724" lane="1" entrytime="00:01:16.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                    <SPLIT distance="75" swimtime="00:00:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="315" swimtime="00:01:21.27" resultid="12647" heatid="14759" lane="2" entrytime="00:01:23.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.54" />
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="75" swimtime="00:01:00.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="359" swimtime="00:01:03.20" resultid="12648" heatid="14790" lane="4" entrytime="00:01:05.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.40" />
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="75" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessio" lastname="Rizzo" birthdate="2010-05-14" gender="M" nation="SUI" license="7982" swrid="5264327" athleteid="12637">
              <RESULTS>
                <RESULT eventid="1081" points="93" swimtime="00:01:46.34" resultid="12638" heatid="14564" lane="2" entrytime="00:01:53.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="115" swimtime="00:01:53.61" resultid="12639" heatid="14622" lane="1" entrytime="00:01:54.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.13" />
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                    <SPLIT distance="75" swimtime="00:01:24.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="109" swimtime="00:01:34.06" resultid="12640" heatid="14673" lane="1" entrytime="00:01:35.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="75" swimtime="00:01:09.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Rossi" birthdate="2004-03-25" gender="M" nation="ITA" license="7999" swrid="5104839" athleteid="12641">
              <RESULTS>
                <RESULT eventid="1111" points="349" swimtime="00:01:07.80" resultid="12642" heatid="14697" lane="1" entrytime="00:01:16.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.75" />
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="75" swimtime="00:00:48.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="364" swimtime="00:01:07.66" resultid="12643" heatid="14727" lane="4" entrytime="00:01:09.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.06" />
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="75" swimtime="00:00:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="470" swimtime="00:00:57.77" resultid="12644" heatid="14794" lane="3" entrytime="00:00:58.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                    <SPLIT distance="75" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliver" lastname="Flüeler" birthdate="2006-03-28" gender="M" nation="SUI" license="8035" swrid="5207277" athleteid="12622">
              <RESULTS>
                <RESULT eventid="1117" points="208" swimtime="00:01:21.48" resultid="12623" heatid="14721" lane="3" entrytime="00:01:26.36">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.43" />
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="75" swimtime="00:01:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="237" swimtime="00:01:29.37" resultid="12624" heatid="14757" lane="2" entrytime="00:01:29.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.95" />
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="75" swimtime="00:01:05.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="339" swimtime="00:01:04.45" resultid="12625" heatid="14789" lane="3" entrytime="00:01:06.63">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.35" />
                    <SPLIT distance="50" swimtime="00:00:30.39" />
                    <SPLIT distance="75" swimtime="00:00:47.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matilda" lastname="Stahl" birthdate="2016-07-07" gender="F" nation="GER" license="42200" swrid="5555306" athleteid="12661">
              <RESULTS>
                <RESULT eventid="1074" status="WDR" swimtime="00:00:00.00" resultid="12662" entrytime="00:01:10.00" />
                <RESULT eventid="1088" status="WDR" swimtime="00:00:00.00" resultid="12663" entrytime="00:01:15.00" />
                <RESULT eventid="1098" status="WDR" swimtime="00:00:00.00" resultid="12664" entrytime="00:01:05.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nico" lastname="Häberli" birthdate="2004-12-18" gender="M" nation="SUI" license="8032" swrid="4892363" athleteid="12626">
              <RESULTS>
                <RESULT eventid="1127" points="466" swimtime="00:01:11.38" resultid="12627" heatid="14761" lane="3" entrytime="00:01:16.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.62" />
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="75" swimtime="00:00:51.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="452" swimtime="00:00:58.55" resultid="12628" heatid="14794" lane="1" entrytime="00:00:58.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.92" />
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                    <SPLIT distance="75" swimtime="00:00:42.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Caligari" birthdate="2014-02-21" gender="F" nation="SUI" license="40905" swrid="5540385" athleteid="12606">
              <RESULTS>
                <RESULT eventid="1074" points="66" swimtime="00:01:03.06" resultid="12607" heatid="14528" lane="2" entrytime="00:01:10.00" />
                <RESULT eventid="1088" points="49" swimtime="00:01:17.67" resultid="12608" heatid="14584" lane="2" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="52" swimtime="00:01:01.42" resultid="12609" heatid="14632" lane="3" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elia" lastname="Stutz" birthdate="2005-01-30" gender="M" nation="SUI" license="11286" swrid="4824776" athleteid="12665">
              <RESULTS>
                <RESULT eventid="1111" points="426" swimtime="00:01:03.50" resultid="12666" heatid="14699" lane="2" entrytime="00:01:04.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.06" />
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="75" swimtime="00:00:46.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="492" swimtime="00:00:56.89" resultid="12667" heatid="14796" lane="4" entrytime="00:00:56.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.65" />
                    <SPLIT distance="50" swimtime="00:00:26.97" />
                    <SPLIT distance="75" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Eigenmann" birthdate="2012-07-05" gender="F" nation="SUI" license="40657" swrid="5555299" athleteid="12618">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="12619" entrytime="00:02:45.00" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="12620" entrytime="00:02:45.00" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="12621" entrytime="00:02:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arsenije" lastname="Arsic" birthdate="2009-05-06" gender="M" nation="SUI" license="7989" swrid="5314251" athleteid="12598">
              <RESULTS>
                <RESULT eventid="1111" points="252" swimtime="00:01:15.64" resultid="12599" heatid="14696" lane="2" entrytime="00:01:22.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.17" />
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="75" swimtime="00:00:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="205" swimtime="00:01:33.80" resultid="12600" heatid="14756" lane="4" entrytime="00:01:35.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.44" />
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                    <SPLIT distance="75" swimtime="00:01:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="248" swimtime="00:01:11.45" resultid="12601" heatid="14787" lane="2" entrytime="00:01:10.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.64" />
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="75" swimtime="00:00:52.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melina" lastname="Zissis" birthdate="2012-02-12" gender="F" nation="SUI" license="8026" swrid="5440453" athleteid="12668">
              <RESULTS>
                <RESULT eventid="1078" points="99" swimtime="00:01:58.63" resultid="12669" heatid="14540" lane="4" entrytime="00:02:05.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="126" swimtime="00:02:04.21" resultid="12670" heatid="14599" lane="1" entrytime="00:02:07.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.48" />
                    <SPLIT distance="50" swimtime="00:00:57.86" />
                    <SPLIT distance="75" swimtime="00:01:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="12671" entrytime="00:01:55.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anne Sophie" lastname="Schweighofer" birthdate="2007-05-24" gender="F" nation="SUI" license="7987" swrid="5264312" athleteid="12657">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 17:11)" eventid="1114" status="DSQ" swimtime="00:01:58.95" resultid="12658" heatid="14703" lane="3" entrytime="00:01:51.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="159" swimtime="00:01:55.09" resultid="12659" heatid="14738" lane="3" entrytime="00:01:56.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.10" />
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                    <SPLIT distance="75" swimtime="00:01:21.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="185" swimtime="00:01:28.06" resultid="12660" heatid="14767" lane="4" entrytime="00:01:25.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.32" />
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rastko" lastname="Arsic" birthdate="2012-06-02" gender="M" nation="SUI" license="32799" swrid="4980890" athleteid="12602">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende 3) (Zeit: 10:25)" eventid="1081" status="DSQ" swimtime="00:02:16.79" resultid="12603" heatid="14560" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.87" />
                    <SPLIT distance="50" swimtime="00:01:01.94" />
                    <SPLIT distance="75" swimtime="00:01:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="57" swimtime="00:02:23.74" resultid="12604" heatid="14617" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.53" />
                    <SPLIT distance="50" swimtime="00:01:07.71" />
                    <SPLIT distance="75" swimtime="00:01:45.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="48" swimtime="00:02:03.63" resultid="12605" heatid="14667" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Palazzoni" birthdate="2007-12-08" gender="F" nation="ITA" license="35808" swrid="5246580" athleteid="12633">
              <RESULTS>
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="12634" entrytime="00:01:42.97" />
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="12635" entrytime="00:01:59.27" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="12636" entrytime="00:01:27.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Diaz" birthdate="2009-11-22" gender="M" nation="SUI" license="19686" swrid="5440436" athleteid="12614">
              <RESULTS>
                <RESULT eventid="1117" points="170" swimtime="00:01:27.22" resultid="12615" heatid="14720" lane="3" entrytime="00:01:31.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.79" />
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="201" swimtime="00:01:34.42" resultid="12616" heatid="14756" lane="1" entrytime="00:01:34.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.71" />
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                    <SPLIT distance="75" swimtime="00:01:08.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="232" swimtime="00:01:13.06" resultid="12617" heatid="14786" lane="2" entrytime="00:01:13.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.36" />
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Schupp" birthdate="2006-11-09" gender="M" nation="SUI" license="8000" swrid="5097306" athleteid="12653">
              <RESULTS>
                <RESULT eventid="1117" points="225" swimtime="00:01:19.44" resultid="12654" heatid="14723" lane="4" entrytime="00:01:22.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.66" />
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="75" swimtime="00:00:58.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...) (Zeit: 18:55)" eventid="1127" status="DSQ" swimtime="00:01:28.63" resultid="12655" heatid="14758" lane="4" entrytime="00:01:29.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.42" />
                    <SPLIT distance="50" swimtime="00:00:41.53" />
                    <SPLIT distance="75" swimtime="00:01:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="267" swimtime="00:01:09.78" resultid="12656" heatid="14789" lane="4" entrytime="00:01:08.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.69" />
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="75" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Loris" lastname="Di Muccio" birthdate="2012-03-23" gender="M" nation="ESP" license="42170" athleteid="12610">
              <RESULTS>
                <RESULT comment="302 - Wand nicht berührt (Wende 2) (Zeit: 10:16)" eventid="1081" status="DSQ" swimtime="00:02:07.12" resultid="12611" heatid="14558" lane="2" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.71" />
                    <SPLIT distance="50" swimtime="00:00:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Zeit: 12:44)" eventid="1095" status="DSQ" swimtime="00:03:19.69" resultid="12612" heatid="14614" lane="3" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:39.89" />
                    <SPLIT distance="50" swimtime="00:01:32.16" />
                    <SPLIT distance="75" swimtime="00:02:24.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="58" swimtime="00:01:55.93" resultid="12613" heatid="14665" lane="1" entrytime="00:04:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.11" />
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                    <SPLIT distance="75" swimtime="00:01:26.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlotta" lastname="Schneider" birthdate="2008-11-11" gender="F" nation="GER" license="7990" swrid="5207266" athleteid="12649">
              <RESULTS>
                <RESULT eventid="1114" points="194" swimtime="00:01:34.80" resultid="12650" heatid="14705" lane="3" entrytime="00:01:33.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.82" />
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="243" swimtime="00:01:39.90" resultid="12651" heatid="14740" lane="3" entrytime="00:01:41.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.07" />
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                    <SPLIT distance="75" swimtime="00:01:12.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="268" swimtime="00:01:17.88" resultid="12652" heatid="14768" lane="2" entrytime="00:01:19.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.50" />
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="75" swimtime="00:00:57.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mila" lastname="Luder" birthdate="2013-03-05" gender="F" nation="SUI" license="32111" swrid="5540389" athleteid="12629">
              <RESULTS>
                <RESULT eventid="1074" status="WDR" swimtime="00:00:00.00" resultid="12630" entrytime="00:00:50.00" />
                <RESULT eventid="1088" status="WDR" swimtime="00:00:00.00" resultid="12631" entrytime="00:00:54.00" />
                <RESULT eventid="1098" status="WDR" swimtime="00:00:00.00" resultid="12632" entrytime="00:00:45.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="453" swimtime="00:01:57.69" resultid="12672" heatid="14736" lane="1" entrytime="00:01:59.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="75" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:03.48" />
                    <SPLIT distance="125" swimtime="00:01:16.20" />
                    <SPLIT distance="150" swimtime="00:01:31.83" />
                    <SPLIT distance="175" swimtime="00:01:44.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12645" number="1" />
                    <RELAYPOSITION athleteid="12626" number="2" />
                    <RELAYPOSITION athleteid="12665" number="3" />
                    <RELAYPOSITION athleteid="12641" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1122" points="283" swimtime="00:02:17.70" resultid="12673" heatid="14735" lane="4" entrytime="00:02:33.20">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="75" swimtime="00:00:54.92" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="125" swimtime="00:01:29.52" />
                    <SPLIT distance="150" swimtime="00:01:47.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12622" number="1" />
                    <RELAYPOSITION athleteid="12653" number="2" />
                    <RELAYPOSITION athleteid="12598" number="3" />
                    <RELAYPOSITION athleteid="12614" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SRSO" nation="SUI" region="RZW" clubid="14325" swrid="87814" name="Swim Regio Solothurn">
          <ATHLETES>
            <ATHLETE firstname="Lea" lastname="Scheidegger" birthdate="2013-05-18" gender="F" nation="SUI" swrid="5564710" athleteid="14420">
              <RESULTS>
                <RESULT eventid="1074" points="101" swimtime="00:00:54.89" resultid="14421" heatid="14530" lane="3" entrytime="00:01:01.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="73" swimtime="00:01:08.06" resultid="14422" heatid="14586" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="95" swimtime="00:00:50.16" resultid="14423" heatid="14635" lane="4" entrytime="00:00:54.92" entrycourse="SCM" />
                <RESULT eventid="1064" points="50" swimtime="00:01:05.98" resultid="14424" heatid="14514" lane="4" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabienne" lastname="Christen" birthdate="2007-04-10" gender="F" nation="SUI" license="102626" swrid="5031991" athleteid="14346">
              <RESULTS>
                <RESULT eventid="1114" points="443" swimtime="00:01:12.00" resultid="14347" heatid="14715" lane="3" entrytime="00:01:10.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.48" />
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="75" swimtime="00:00:53.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="472" swimtime="00:01:04.53" resultid="14348" heatid="14777" lane="2" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.67" />
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="75" swimtime="00:00:47.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Selina" lastname="Rickli" birthdate="2008-07-23" gender="F" nation="SUI" license="108728" swrid="5151072" athleteid="14411">
              <RESULTS>
                <RESULT eventid="1108" points="197" swimtime="00:01:33.82" resultid="14412" heatid="14685" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.76" />
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                    <SPLIT distance="75" swimtime="00:01:09.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="228" swimtime="00:01:29.73" resultid="14413" heatid="14708" lane="3" entrytime="00:01:24.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.37" />
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="75" swimtime="00:01:07.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="215" swimtime="00:01:44.00" resultid="14414" heatid="14741" lane="1" entrytime="00:01:39.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.33" />
                    <SPLIT distance="50" swimtime="00:00:51.38" />
                    <SPLIT distance="75" swimtime="00:01:17.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="303" swimtime="00:01:14.77" resultid="14415" heatid="14771" lane="3" entrytime="00:01:12.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.34" />
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="75" swimtime="00:00:56.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noée" lastname="Lombardi" birthdate="2014-07-23" gender="F" nation="SUI" license="38628" swrid="5497470" athleteid="14395">
              <RESULTS>
                <RESULT eventid="1074" points="78" swimtime="00:00:59.75" resultid="14396" heatid="14531" lane="1" entrytime="00:00:59.96" entrycourse="LCM" />
                <RESULT eventid="1098" points="73" swimtime="00:00:54.64" resultid="14397" heatid="14635" lane="3" entrytime="00:00:53.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Zeit: 11:54)" eventid="1088" status="DSQ" swimtime="00:01:11.42" resultid="14398" heatid="14588" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matej" lastname="Niznik" birthdate="2009-01-20" gender="M" nation="SVK" license="7067" swrid="5398274" athleteid="14406">
              <RESULTS>
                <RESULT eventid="1111" points="255" swimtime="00:01:15.29" resultid="14407" heatid="14697" lane="4" entrytime="00:01:22.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.30" />
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="75" swimtime="00:00:55.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="235" swimtime="00:01:18.30" resultid="14408" heatid="14721" lane="1" entrytime="00:01:29.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.74" />
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="75" swimtime="00:00:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="316" swimtime="00:01:21.20" resultid="14409" heatid="14760" lane="1" entrytime="00:01:22.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.44" />
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="75" swimtime="00:00:59.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="318" swimtime="00:01:05.84" resultid="14410" heatid="14789" lane="2" entrytime="00:01:05.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.13" />
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="75" swimtime="00:00:49.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fiona Sophia" lastname="Eterno" birthdate="2010-02-09" gender="F" nation="SUI" license="27326" swrid="5464162" athleteid="14360">
              <RESULTS>
                <RESULT eventid="1078" points="191" swimtime="00:01:35.31" resultid="14361" heatid="14546" lane="3" entrytime="00:01:44.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="140" swimtime="00:02:00.01" resultid="14362" heatid="14600" lane="1" entrytime="00:02:04.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.33" />
                    <SPLIT distance="50" swimtime="00:00:54.83" />
                    <SPLIT distance="75" swimtime="00:01:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="178" swimtime="00:01:29.25" resultid="14363" heatid="14648" lane="4" entrytime="00:01:41.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.10" />
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="75" swimtime="00:01:05.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Schor" birthdate="2012-10-13" gender="M" nation="SUI" swrid="5231088" athleteid="14425">
              <RESULTS>
                <RESULT eventid="1081" points="63" swimtime="00:02:00.84" resultid="14426" heatid="14567" lane="4" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.71" />
                    <SPLIT distance="50" swimtime="00:00:57.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="58" swimtime="00:02:22.92" resultid="14427" heatid="14617" lane="1" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:32.19" />
                    <SPLIT distance="50" swimtime="00:01:09.09" />
                    <SPLIT distance="75" swimtime="00:01:47.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="61" swimtime="00:01:53.97" resultid="14428" heatid="14671" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Seraina" lastname="Häfliger" birthdate="2012-08-14" gender="F" nation="SUI" license="19309" swrid="5464167" athleteid="14375">
              <RESULTS>
                <RESULT eventid="1078" points="152" swimtime="00:01:42.71" resultid="14376" heatid="14545" lane="3" entrytime="00:01:45.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.19" />
                    <SPLIT distance="75" swimtime="00:01:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="111" swimtime="00:02:09.69" resultid="14377" heatid="14598" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.06" />
                    <SPLIT distance="50" swimtime="00:00:59.27" />
                    <SPLIT distance="75" swimtime="00:01:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="145" swimtime="00:01:35.56" resultid="14378" heatid="14647" lane="2" entrytime="00:01:43.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.21" />
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                    <SPLIT distance="75" swimtime="00:01:12.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valerie" lastname="Bur" birthdate="2013-09-09" gender="F" nation="SUI" license="32336" swrid="5484580" athleteid="14342">
              <RESULTS>
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="14343" heatid="14529" lane="1" entrytime="00:01:07.03" entrycourse="SCM" />
                <RESULT eventid="1088" status="DNS" swimtime="00:00:00.00" resultid="14344" heatid="14585" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="14345" heatid="14633" lane="2" entrytime="00:00:58.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melanie" lastname="Christen" birthdate="2011-10-04" gender="F" nation="SUI" license="116469" swrid="5263509" athleteid="14349">
              <RESULTS>
                <RESULT eventid="1068" points="116" swimtime="00:01:51.75" resultid="14350" heatid="14518" lane="2" entrytime="00:01:50.10">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.39" />
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="75" swimtime="00:01:20.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="176" swimtime="00:01:51.07" resultid="14351" heatid="14606" lane="3" entrytime="00:01:42.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.89" />
                    <SPLIT distance="50" swimtime="00:00:52.25" />
                    <SPLIT distance="75" swimtime="00:01:21.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="193" swimtime="00:01:26.85" resultid="14352" heatid="14653" lane="3" entrytime="00:01:27.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.93" />
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="75" swimtime="00:01:04.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Wyss" birthdate="2012-03-18" gender="M" nation="SUI" license="7087" swrid="5411009" athleteid="14447">
              <RESULTS>
                <RESULT eventid="1081" points="113" swimtime="00:01:39.68" resultid="14448" heatid="14569" lane="1" entrytime="00:01:40.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.34" />
                    <SPLIT distance="50" swimtime="00:00:48.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="117" swimtime="00:01:53.14" resultid="14449" heatid="14618" lane="2" entrytime="00:02:09.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.73" />
                    <SPLIT distance="50" swimtime="00:00:55.00" />
                    <SPLIT distance="75" swimtime="00:01:24.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="123" swimtime="00:01:30.30" resultid="14450" heatid="14671" lane="1" entrytime="00:01:40.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.13" />
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="75" swimtime="00:01:09.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefanie" lastname="Christen" birthdate="2009-01-30" gender="F" nation="SUI" license="107842" swrid="5151069" athleteid="14353">
              <RESULTS>
                <RESULT eventid="1108" points="240" swimtime="00:01:27.87" resultid="14354" heatid="14685" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.61" />
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="75" swimtime="00:01:02.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="336" swimtime="00:01:18.94" resultid="14355" heatid="14709" lane="3" entrytime="00:01:21.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                    <SPLIT distance="75" swimtime="00:00:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="400" swimtime="00:01:08.18" resultid="14356" heatid="14774" lane="2" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.31" />
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="75" swimtime="00:00:50.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gaetano" lastname="Furrer" birthdate="2012-09-13" gender="M" nation="SUI" license="19166" swrid="5464164" athleteid="14364">
              <RESULTS>
                <RESULT eventid="1081" points="113" swimtime="00:01:39.96" resultid="14365" heatid="14564" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.76" />
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="84" swimtime="00:02:06.27" resultid="14366" heatid="14618" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.23" />
                    <SPLIT distance="50" swimtime="00:01:02.04" />
                    <SPLIT distance="75" swimtime="00:01:34.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="108" swimtime="00:01:34.15" resultid="14367" heatid="14669" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.85" />
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="75" swimtime="00:01:10.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elin" lastname="Gerber" birthdate="2011-03-13" gender="F" nation="SUI" license="27005" swrid="5509051" athleteid="14368">
              <RESULTS>
                <RESULT eventid="1078" points="119" swimtime="00:01:51.33" resultid="14369" heatid="14544" lane="4" entrytime="00:01:49.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.93" />
                    <SPLIT distance="50" swimtime="00:00:53.55" />
                    <SPLIT distance="75" swimtime="00:01:22.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="133" swimtime="00:01:38.29" resultid="14370" heatid="14648" lane="2" entrytime="00:01:39.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.29" />
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adina" lastname="Schütz" birthdate="2010-05-26" gender="F" nation="SUI" license="37863" swrid="5509054" athleteid="14429">
              <RESULTS>
                <RESULT eventid="1078" points="167" swimtime="00:01:39.49" resultid="14430" heatid="14544" lane="3" entrytime="00:01:48.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="257" swimtime="00:01:37.99" resultid="14431" heatid="14605" lane="2" entrytime="00:01:44.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.35" />
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                    <SPLIT distance="75" swimtime="00:01:11.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="205" swimtime="00:01:25.17" resultid="14432" heatid="14650" lane="1" entrytime="00:01:38.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="75" swimtime="00:01:02.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lenny" lastname="Steiner" birthdate="2012-03-09" gender="M" nation="SUI" license="28648" swrid="5464191" athleteid="14433">
              <RESULTS>
                <RESULT eventid="1081" points="93" swimtime="00:01:46.34" resultid="14434" heatid="14563" lane="2" entrytime="00:01:57.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="128" swimtime="00:01:49.65" resultid="14435" heatid="14623" lane="1" entrytime="00:01:53.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.72" />
                    <SPLIT distance="50" swimtime="00:00:52.87" />
                    <SPLIT distance="75" swimtime="00:01:20.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="90" swimtime="00:01:40.10" resultid="14436" heatid="14668" lane="1" entrytime="00:01:55.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.13" />
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                    <SPLIT distance="75" swimtime="00:01:13.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Kurth" birthdate="2013-06-02" gender="F" nation="SUI" license="19263" swrid="5464176" athleteid="14383">
              <RESULTS>
                <RESULT comment="505 - Wechselbeinschlag während des Schwimmens (Zeit: 8:43)" eventid="1064" status="DSQ" swimtime="00:01:02.93" resultid="14384" heatid="14514" lane="1" entrytime="00:00:59.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 9:19)" eventid="1074" status="DSQ" swimtime="00:00:54.08" resultid="14385" heatid="14532" lane="3" entrytime="00:00:54.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="117" swimtime="00:00:46.82" resultid="14386" heatid="14636" lane="1" entrytime="00:00:47.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="107" swimtime="00:01:00.00" resultid="14387" heatid="14588" lane="1" entrytime="00:01:02.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabella" lastname="Elias" birthdate="2011-05-05" gender="F" nation="HUN" license="19004" swrid="5540421" athleteid="14357">
              <RESULTS>
                <RESULT eventid="1102" points="105" swimtime="00:01:46.38" resultid="14358" heatid="14647" lane="4" entrytime="00:01:47.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.84" />
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                    <SPLIT distance="75" swimtime="00:01:18.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="75" swimtime="00:02:10.09" resultid="14359" heatid="14539" lane="2" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.76" />
                    <SPLIT distance="50" swimtime="00:01:01.28" />
                    <SPLIT distance="75" swimtime="00:01:36.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Würgler" birthdate="2009-06-29" gender="F" nation="SUI" license="7116" swrid="5395766" athleteid="14442">
              <RESULTS>
                <RESULT eventid="1114" points="224" swimtime="00:01:30.31" resultid="14443" heatid="14706" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="404" swimtime="00:01:24.30" resultid="14444" heatid="14746" lane="2" entrytime="00:01:27.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.35" />
                    <SPLIT distance="50" swimtime="00:00:39.52" />
                    <SPLIT distance="75" swimtime="00:01:01.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="338" swimtime="00:01:12.11" resultid="14445" heatid="14772" lane="1" entrytime="00:01:11.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.96" />
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="75" swimtime="00:00:54.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1108" points="219" swimtime="00:01:30.59" resultid="14446" heatid="14685" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.49" />
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="75" swimtime="00:01:04.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Céline" lastname="Torre" birthdate="2013-04-08" gender="F" nation="SUI" license="19172" swrid="5464194" athleteid="14437">
              <RESULTS>
                <RESULT eventid="1074" points="83" swimtime="00:00:58.56" resultid="14438" heatid="14530" lane="1" entrytime="00:01:01.76" entrycourse="LCM" />
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...) (Zeit: 11:58)" eventid="1088" status="DSQ" swimtime="00:01:06.30" resultid="14439" heatid="14587" lane="4" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="76" swimtime="00:00:53.96" resultid="14440" heatid="14634" lane="3" entrytime="00:00:56.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="52" swimtime="00:01:05.05" resultid="14441" heatid="14513" lane="2" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia Sarai" lastname="Günther" birthdate="2011-11-29" gender="F" nation="SUI" license="121779" swrid="5411028" athleteid="14371">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="14372" entrytime="00:01:52.35" entrycourse="SCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="14373" entrytime="00:01:50.78" entrycourse="SCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="14374" entrytime="00:01:40.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lars" lastname="Lyszczynski" birthdate="2011-06-15" gender="M" nation="SUI" license="19261" swrid="5540422" athleteid="14399">
              <RESULTS>
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="14400" entrytime="00:02:10.00" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="14401" entrytime="00:01:42.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nia Mara" lastname="Lemp" birthdate="2011-05-19" gender="F" nation="SUI" license="19118" swrid="5467814" athleteid="14391">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 10:30)" eventid="1078" status="DSQ" swimtime="00:01:48.08" resultid="14392" heatid="14541" lane="4" entrytime="00:02:03.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.79" />
                    <SPLIT distance="50" swimtime="00:00:50.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="114" swimtime="00:02:08.32" resultid="14393" heatid="14597" lane="4" entrytime="00:02:16.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.76" />
                    <SPLIT distance="50" swimtime="00:01:01.34" />
                    <SPLIT distance="75" swimtime="00:01:34.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="123" swimtime="00:01:40.97" resultid="14394" heatid="14646" lane="3" entrytime="00:01:50.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.04" />
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                    <SPLIT distance="75" swimtime="00:01:15.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lean" lastname="Müller" birthdate="2013-06-28" gender="M" nation="SUI" license="28040" swrid="5523508" athleteid="14402">
              <RESULTS>
                <RESULT eventid="1076" points="60" swimtime="00:00:56.51" resultid="14403" heatid="14536" lane="2" entrytime="00:00:57.57" entrycourse="SCM" />
                <RESULT eventid="1090" points="79" swimtime="00:00:58.70" resultid="14404" heatid="14594" lane="4" entrytime="00:00:59.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="62" swimtime="00:00:50.88" resultid="14405" heatid="14639" lane="2" entrytime="00:00:52.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pascal" lastname="Zollinger" birthdate="2001-03-16" gender="M" nation="SUI" license="46474" swrid="4879834" athleteid="14451">
              <RESULTS>
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="14452" entrytime="00:01:05.61" entrycourse="SCM" />
                <RESULT eventid="1117" points="402" swimtime="00:01:05.44" resultid="14453" heatid="14727" lane="2" entrytime="00:01:08.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.03" />
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="75" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" status="WDR" swimtime="00:00:00.00" resultid="14454" entrytime="00:01:13.57" entrycourse="SCM" />
                <RESULT eventid="1133" points="568" swimtime="00:00:54.25" resultid="14455" heatid="14796" lane="2" entrytime="00:00:54.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.41" />
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                    <SPLIT distance="75" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="382" swimtime="00:00:30.60" resultid="14852" heatid="14802" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6683" points="459" swimtime="00:00:32.73" resultid="14867" heatid="14804" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mailey Sue" lastname="Bruns" birthdate="2011-09-12" gender="F" nation="GER" license="120076" swrid="5329307" athleteid="14338">
              <RESULTS>
                <RESULT eventid="1078" points="324" swimtime="00:01:19.87" resultid="14339" heatid="14554" lane="4" entrytime="00:01:19.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.04" />
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="75" swimtime="00:00:58.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="257" swimtime="00:01:38.02" resultid="14340" heatid="14607" lane="2" entrytime="00:01:38.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.60" />
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                    <SPLIT distance="75" swimtime="00:01:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="389" swimtime="00:01:08.80" resultid="14341" heatid="14661" lane="4" entrytime="00:01:10.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.25" />
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="75" swimtime="00:00:50.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucia" lastname="Rinaldi" birthdate="2009-12-21" gender="F" nation="SUI" license="40440" swrid="5521571" athleteid="14416">
              <RESULTS>
                <RESULT eventid="1114" points="113" swimtime="00:01:53.39" resultid="14417" heatid="14703" lane="1" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="130" swimtime="00:02:02.97" resultid="14418" heatid="14738" lane="1" entrytime="00:02:02.78">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.31" />
                    <SPLIT distance="50" swimtime="00:00:58.08" />
                    <SPLIT distance="75" swimtime="00:01:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="140" swimtime="00:01:36.55" resultid="14419" heatid="14765" lane="3" entrytime="00:01:36.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.09" />
                    <SPLIT distance="50" swimtime="00:00:45.02" />
                    <SPLIT distance="75" swimtime="00:01:12.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mira" lastname="Leibundgut" birthdate="2008-09-20" gender="F" nation="SUI" license="107744" swrid="5133787" athleteid="14388">
              <RESULTS>
                <RESULT eventid="1124" points="333" swimtime="00:01:29.93" resultid="14389" heatid="14747" lane="1" entrytime="00:01:26.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.32" />
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                    <SPLIT distance="75" swimtime="00:01:05.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="403" swimtime="00:01:08.01" resultid="14390" heatid="14775" lane="4" entrytime="00:01:08.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caroline Mathilde" lastname="Bang" birthdate="2006-10-15" gender="F" nation="DEN" license="116476" swrid="5057737" athleteid="14331">
              <RESULTS>
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="14332" entrytime="00:01:01.26" entrycourse="SCM" />
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="14333" entrytime="00:01:10.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Levi" lastname="Berger" birthdate="2013-04-03" gender="M" nation="SUI" license="19071" swrid="5464156" athleteid="14334">
              <RESULTS>
                <RESULT eventid="1076" points="57" swimtime="00:00:57.43" resultid="14335" heatid="14535" lane="3" entrytime="00:01:01.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="60" swimtime="00:00:51.48" resultid="14336" heatid="14640" lane="2" entrytime="00:00:48.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="26" swimtime="00:01:25.22" resultid="14337" heatid="14592" lane="1" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:35.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Naira" lastname="Kägi" birthdate="2011-08-05" gender="F" nation="SUI" license="121390" swrid="5353510" athleteid="14379">
              <RESULTS>
                <RESULT eventid="1068" points="128" swimtime="00:01:48.29" resultid="14380" heatid="14518" lane="1" entrytime="00:01:56.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.54" />
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                    <SPLIT distance="75" swimtime="00:01:19.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="217" swimtime="00:01:31.32" resultid="14381" heatid="14551" lane="1" entrytime="00:01:35.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.36" />
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="75" swimtime="00:01:08.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="225" swimtime="00:01:22.58" resultid="14382" heatid="14654" lane="1" entrytime="00:01:26.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.06" />
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="75" swimtime="00:01:01.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eliott" lastname="André" birthdate="2007-10-13" gender="M" nation="SUI" license="19313" swrid="5467808" athleteid="14326">
              <RESULTS>
                <RESULT eventid="1111" points="331" swimtime="00:01:09.02" resultid="14327" heatid="14698" lane="4" entrytime="00:01:10.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.20" />
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="75" swimtime="00:00:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="351" swimtime="00:01:08.48" resultid="14328" heatid="14726" lane="1" entrytime="00:01:11.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.45" />
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                    <SPLIT distance="75" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="303" swimtime="00:01:22.35" resultid="14329" heatid="14758" lane="2" entrytime="00:01:25.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.76" />
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="75" swimtime="00:01:00.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="349" swimtime="00:01:03.77" resultid="14330" heatid="14791" lane="4" entrytime="00:01:04.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.48" />
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="75" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 11:33)" eventid="1086" status="DSQ" swimtime="00:02:55.29" resultid="14456" heatid="14582" lane="1" entrytime="00:02:53.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.10" />
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="75" swimtime="00:01:01.01" />
                    <SPLIT distance="100" swimtime="00:01:23.74" />
                    <SPLIT distance="125" swimtime="00:01:42.66" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                    <SPLIT distance="175" swimtime="00:02:28.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14447" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="14364" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="14433" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="14425" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="248" swimtime="00:02:27.11" resultid="14457" heatid="14580" lane="1" entrytime="00:02:30.57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.84" />
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="75" swimtime="00:00:49.29" />
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                    <SPLIT distance="125" swimtime="00:01:29.56" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                    <SPLIT distance="175" swimtime="00:02:07.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14338" number="1" />
                    <RELAYPOSITION athleteid="14379" number="2" />
                    <RELAYPOSITION athleteid="14375" number="3" />
                    <RELAYPOSITION athleteid="14349" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="425" swimtime="00:02:16.08" resultid="14458" heatid="14733" lane="1" entrytime="00:02:11.52">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.60" />
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="75" swimtime="00:00:51.01" />
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                    <SPLIT distance="125" swimtime="00:01:27.20" />
                    <SPLIT distance="150" swimtime="00:01:45.52" />
                    <SPLIT distance="175" swimtime="00:02:00.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14346" number="1" />
                    <RELAYPOSITION athleteid="14442" number="2" />
                    <RELAYPOSITION athleteid="14388" number="3" />
                    <RELAYPOSITION athleteid="14353" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1084" points="182" swimtime="00:02:42.94" resultid="14459" heatid="14578" lane="1" entrytime="00:02:54.03">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.52" />
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="75" swimtime="00:00:57.83" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="125" swimtime="00:01:39.07" />
                    <SPLIT distance="150" swimtime="00:01:58.92" />
                    <SPLIT distance="175" swimtime="00:02:19.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14429" number="1" />
                    <RELAYPOSITION athleteid="14391" number="2" />
                    <RELAYPOSITION athleteid="14360" number="3" />
                    <RELAYPOSITION athleteid="14368" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer 4) (Zeit: 11:16)" eventid="1084" status="DSQ" swimtime="00:03:24.15" resultid="14460" heatid="14576" lane="2" entrytime="00:03:31.57">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.41" />
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                    <SPLIT distance="75" swimtime="00:01:13.86" />
                    <SPLIT distance="100" swimtime="00:01:43.48" />
                    <SPLIT distance="125" swimtime="00:02:54.62" />
                    <SPLIT distance="150" swimtime="00:02:33.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14383" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="14395" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="14420" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="14437" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ALL" nation="SUI" region="RZW" clubid="13363" swrid="65684" name="Schwimmclub Allschwil">
          <ATHLETES>
            <ATHLETE firstname="David" lastname="Beshai" birthdate="2010-10-19" gender="M" nation="SUI" license="33046" swrid="5564693" athleteid="13364">
              <RESULTS>
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="13365" entrytime="00:01:42.77" />
                <RESULT eventid="1095" status="WDR" swimtime="00:00:00.00" resultid="13366" entrytime="00:01:55.00" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="13367" entrytime="00:01:40.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Di Ciancia Ferreira" birthdate="2013-05-19" gender="F" nation="SUI" license="33588" swrid="5564696" athleteid="13375">
              <RESULTS>
                <RESULT eventid="1074" points="94" swimtime="00:00:56.29" resultid="13376" heatid="14530" lane="2" entrytime="00:01:00.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="68" swimtime="00:01:09.90" resultid="13377" heatid="14587" lane="1" entrytime="00:01:09.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="78" swimtime="00:00:53.65" resultid="13378" heatid="14634" lane="2" entrytime="00:00:56.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Chloé" lastname="Duréault" birthdate="2008-02-28" gender="F" nation="SUI" license="37631" swrid="5281922" athleteid="13379">
              <RESULTS>
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="13380" entrytime="00:01:22.71" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="13381" entrytime="00:01:10.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nils" lastname="Schütz" birthdate="2010-11-03" gender="M" nation="SUI" license="32580" swrid="5467817" athleteid="13386">
              <RESULTS>
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="13387" entrytime="00:01:44.05" entrycourse="SCM" />
                <RESULT eventid="1095" status="WDR" swimtime="00:00:00.00" resultid="13388" entrytime="00:01:49.59" entrycourse="SCM" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="13389" entrytime="00:01:37.04" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliver" lastname="Story" birthdate="2007-07-03" gender="M" nation="SUI" license="6592" swrid="5395754" athleteid="13390">
              <RESULTS>
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="13391" entrytime="00:01:19.35" entrycourse="SCM" />
                <RESULT eventid="1133" status="WDR" swimtime="00:00:00.00" resultid="13392" entrytime="00:01:08.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alvaro" lastname="Cancela" birthdate="2009-02-21" gender="M" nation="SUI" license="6375" swrid="5255603" athleteid="13372">
              <RESULTS>
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="13373" entrytime="00:01:20.33" entrycourse="SCM" />
                <RESULT eventid="1133" status="WDR" swimtime="00:00:00.00" resultid="13374" entrytime="00:01:05.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matti" lastname="Brigger" birthdate="2010-06-28" gender="M" nation="SUI" license="32346" swrid="4000990" athleteid="13368">
              <RESULTS>
                <RESULT eventid="1081" points="117" swimtime="00:01:38.59" resultid="13369" heatid="14568" lane="2" entrytime="00:01:42.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.37" />
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="75" swimtime="00:01:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="111" swimtime="00:01:55.08" resultid="13370" heatid="14625" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.66" />
                    <SPLIT distance="50" swimtime="00:00:53.74" />
                    <SPLIT distance="75" swimtime="00:01:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="120" swimtime="00:01:30.90" resultid="13371" heatid="14674" lane="3" entrytime="00:01:33.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.96" />
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="75" swimtime="00:01:08.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amélie" lastname="Grillon" birthdate="2009-04-28" gender="F" nation="SUI" license="6376" swrid="5398284" athleteid="13382">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="13383" entrytime="00:01:26.56" entrycourse="SCM" />
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="13384" entrytime="00:01:25.56" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="13385" entrytime="00:01:09.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="WAED" nation="SUI" region="RZO" clubid="12955" swrid="65647" name="Schwimmverein Wädenswil">
          <ATHLETES>
            <ATHLETE firstname="Tara" lastname="Alberts" birthdate="2013-09-12" gender="F" nation="SUI" license="40644" swrid="5508979" athleteid="12956">
              <RESULTS>
                <RESULT eventid="1064" points="136" swimtime="00:00:47.39" resultid="12957" heatid="14515" lane="4" entrytime="00:00:52.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="132" swimtime="00:00:50.25" resultid="12958" heatid="14532" lane="2" entrytime="00:00:51.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="145" swimtime="00:00:54.30" resultid="12959" heatid="14588" lane="3" entrytime="00:00:59.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="156" swimtime="00:00:42.52" resultid="12960" heatid="14636" lane="2" entrytime="00:00:44.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luciano" lastname="Kick Bedoya" birthdate="2011-09-29" gender="M" nation="GER" license="21194" swrid="5458198" athleteid="13046">
              <RESULTS>
                <RESULT eventid="1081" points="66" swimtime="00:01:59.25" resultid="13047" heatid="14560" lane="2" entrytime="00:02:06.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.87" />
                    <SPLIT distance="50" swimtime="00:00:55.35" />
                    <SPLIT distance="75" swimtime="00:01:27.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="60" swimtime="00:02:21.29" resultid="13048" heatid="14620" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.88" />
                    <SPLIT distance="50" swimtime="00:01:05.01" />
                    <SPLIT distance="75" swimtime="00:01:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="54" swimtime="00:01:58.60" resultid="13049" heatid="14669" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.37" />
                    <SPLIT distance="50" swimtime="00:00:53.94" />
                    <SPLIT distance="75" swimtime="00:01:26.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tymofii" firstname.en="Timothy" lastname="Kozhanov" birthdate="2010-09-16" gender="M" nation="UKR" license="43093" athleteid="13050">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende 3) (Zeit: 10:46)" eventid="1081" status="DSQ" swimtime="00:01:43.57" resultid="13051" heatid="14570" lane="4" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                    <SPLIT distance="75" swimtime="00:01:17.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Nicht mit beiden Händen gleichzeitig angeschlagen (Ziel) (Zeit: 13:24)" eventid="1095" status="DSQ" swimtime="00:02:00.08" resultid="13052" heatid="14626" lane="4" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.45" />
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                    <SPLIT distance="75" swimtime="00:01:27.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="124" swimtime="00:01:30.11" resultid="13053" heatid="14673" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.78" />
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="75" swimtime="00:01:05.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martin" lastname="Dickhoff" birthdate="2006-04-07" gender="M" nation="FRA" license="5725" swrid="5209648" athleteid="12996">
              <RESULTS>
                <RESULT eventid="1117" points="260" swimtime="00:01:15.68" resultid="12997" heatid="14724" lane="3" entrytime="00:01:15.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.59" />
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="241" swimtime="00:01:28.89" resultid="12998" heatid="14756" lane="2" entrytime="00:01:34.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.34" />
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                    <SPLIT distance="75" swimtime="00:01:04.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="319" swimtime="00:01:05.71" resultid="12999" heatid="14791" lane="1" entrytime="00:01:03.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.31" />
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                    <SPLIT distance="75" swimtime="00:00:48.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wanglen" lastname="Mendro" birthdate="2010-05-27" gender="M" nation="SUI" license="5763" swrid="4596908" athleteid="13062">
              <RESULTS>
                <RESULT eventid="1081" points="84" status="DNS" swimtime="00:01:50.04" resultid="13063" heatid="14565" lane="3" entrytime="00:01:49.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="13064" heatid="14622" lane="2" entrytime="00:01:54.06" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="13065" heatid="14677" lane="2" entrytime="00:01:26.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Graser" birthdate="2009-02-01" gender="F" nation="GER" license="5717" swrid="4607405" athleteid="13000">
              <RESULTS>
                <RESULT eventid="1114" points="270" swimtime="00:01:24.84" resultid="13001" heatid="14707" lane="2" entrytime="00:01:25.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.82" />
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="339" swimtime="00:01:29.40" resultid="13002" heatid="14746" lane="4" entrytime="00:01:29.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.22" />
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="75" swimtime="00:01:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="327" swimtime="00:01:12.92" resultid="13003" heatid="14770" lane="1" entrytime="00:01:14.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.73" />
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="75" swimtime="00:00:54.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Evi" lastname="Chambers" birthdate="2009-04-18" gender="F" nation="SUI" license="5685" swrid="4415887" athleteid="12982">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="12983" heatid="14684" lane="3" entrytime="00:01:40.00" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="12984" heatid="14707" lane="1" entrytime="00:01:27.82" entrycourse="SCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="12985" heatid="14743" lane="4" entrytime="00:01:33.63" entrycourse="SCM" />
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="12986" heatid="14770" lane="4" entrytime="00:01:15.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anina" lastname="Werlen" birthdate="2008-04-25" gender="F" nation="SUI" license="5662" swrid="4941067" athleteid="13142">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende 2) (Zeit: 17:26)" eventid="1114" status="DSQ" swimtime="00:01:21.27" resultid="13143" heatid="14709" lane="1" entrytime="00:01:22.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="75" swimtime="00:01:00.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="292" swimtime="00:01:33.90" resultid="13144" heatid="14743" lane="2" entrytime="00:01:32.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.17" />
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="75" swimtime="00:01:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="324" swimtime="00:01:13.09" resultid="13145" heatid="14770" lane="2" entrytime="00:01:13.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.95" />
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="75" swimtime="00:00:54.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leona" lastname="Papp" birthdate="2009-07-09" gender="F" nation="HUN" license="5707" swrid="5351841" athleteid="13083">
              <RESULTS>
                <RESULT eventid="1108" points="418" swimtime="00:01:12.98" resultid="13084" heatid="14690" lane="4" entrytime="00:01:15.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.60" />
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="75" swimtime="00:00:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="304" swimtime="00:01:32.74" resultid="13085" heatid="14744" lane="3" entrytime="00:01:31.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.45" />
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                    <SPLIT distance="75" swimtime="00:01:08.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="557" swimtime="00:01:06.71" resultid="13086" heatid="14716" lane="1" entrytime="00:01:05.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.40" />
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                    <SPLIT distance="75" swimtime="00:00:49.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="518" swimtime="00:01:02.55" resultid="13087" heatid="14780" lane="3" entrytime="00:01:01.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.08" />
                    <SPLIT distance="50" swimtime="00:00:29.89" />
                    <SPLIT distance="75" swimtime="00:00:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="543" swimtime="00:00:31.37" resultid="14844" heatid="14801" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanni" lastname="Mendola" birthdate="2008-08-28" gender="M" nation="ITA" license="43022" swrid="5178015" athleteid="13058">
              <RESULTS>
                <RESULT eventid="1117" points="268" swimtime="00:01:14.88" resultid="13059" heatid="14723" lane="2" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.89" />
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="75" swimtime="00:00:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="212" swimtime="00:01:32.70" resultid="13060" heatid="14757" lane="4" entrytime="00:01:31.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.11" />
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="75" swimtime="00:01:07.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="279" swimtime="00:01:08.76" resultid="13061" heatid="14788" lane="4" entrytime="00:01:10.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.62" />
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="75" swimtime="00:00:51.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrea" lastname="D&apos; Ignazio" birthdate="2007-07-09" gender="M" nation="ITA" license="5661" swrid="5266505" athleteid="12991">
              <RESULTS>
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="12992" heatid="14698" lane="3" entrytime="00:01:09.52" entrycourse="SCM" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="12993" heatid="14725" lane="4" entrytime="00:01:14.58" entrycourse="SCM" />
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="12994" heatid="14761" lane="4" entrytime="00:01:17.53" entrycourse="SCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="12995" heatid="14793" lane="4" entrytime="00:01:00.18" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erik" lastname="Tattersall" birthdate="2011-07-12" gender="M" nation="SUI" license="5683" swrid="5351137" athleteid="13133">
              <RESULTS>
                <RESULT eventid="1071" status="WDR" swimtime="00:00:00.00" resultid="13134" entrytime="00:01:50.00" />
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="13135" entrytime="00:01:50.88" entrycourse="LCM" />
                <RESULT eventid="1095" status="WDR" swimtime="00:00:00.00" resultid="13136" entrytime="00:01:48.19" entrycourse="LCM" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="13137" entrytime="00:01:33.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celine" lastname="Hutter" birthdate="2011-01-04" gender="F" nation="SUI" license="5670" swrid="5351135" athleteid="13012">
              <RESULTS>
                <RESULT eventid="1078" points="203" swimtime="00:01:33.35" resultid="13013" heatid="14549" lane="1" entrytime="00:01:37.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.49" />
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="75" swimtime="00:01:09.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="233" swimtime="00:01:41.31" resultid="13014" heatid="14608" lane="2" entrytime="00:01:35.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.12" />
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                    <SPLIT distance="75" swimtime="00:01:13.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="239" swimtime="00:01:20.94" resultid="13015" heatid="14656" lane="4" entrytime="00:01:24.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.99" />
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Papp" birthdate="2013-05-10" gender="F" nation="HUN" license="32023" swrid="5458213" athleteid="13078">
              <RESULTS>
                <RESULT eventid="1064" points="197" swimtime="00:00:41.86" resultid="13079" heatid="14515" lane="3" entrytime="00:00:49.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="231" swimtime="00:00:41.67" resultid="13080" heatid="14533" lane="2" entrytime="00:00:43.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="245" swimtime="00:00:45.59" resultid="13081" heatid="14589" lane="2" entrytime="00:00:44.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="243" swimtime="00:00:36.71" resultid="13082" heatid="14637" lane="2" entrytime="00:00:35.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Frederic" lastname="Reiter" birthdate="2008-12-19" gender="M" nation="SUI" license="5689" swrid="5242698" athleteid="13097">
              <RESULTS>
                <RESULT eventid="1117" points="201" swimtime="00:01:22.48" resultid="13098" heatid="14723" lane="1" entrytime="00:01:21.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.54" />
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="75" swimtime="00:01:01.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="250" swimtime="00:01:11.33" resultid="13099" heatid="14787" lane="1" entrytime="00:01:11.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.07" />
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                    <SPLIT distance="75" swimtime="00:00:53.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julienne" lastname="Hutter" birthdate="2013-08-03" gender="F" nation="SUI" license="21191" swrid="5440821" athleteid="13016">
              <RESULTS>
                <RESULT eventid="1064" points="147" swimtime="00:00:46.12" resultid="13017" heatid="14515" lane="2" entrytime="00:00:47.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="178" swimtime="00:00:45.46" resultid="13018" heatid="14533" lane="3" entrytime="00:00:45.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="167" swimtime="00:00:51.82" resultid="13019" heatid="14589" lane="1" entrytime="00:00:53.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="270" swimtime="00:00:35.44" resultid="13020" heatid="14637" lane="3" entrytime="00:00:38.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Zellweger" birthdate="2012-09-11" gender="M" nation="SUI" license="32032" swrid="5458232" athleteid="13158">
              <RESULTS>
                <RESULT eventid="1081" points="99" swimtime="00:01:44.17" resultid="13159" heatid="14561" lane="1" entrytime="00:02:06.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.88" />
                    <SPLIT distance="50" swimtime="00:00:52.26" />
                    <SPLIT distance="75" swimtime="00:01:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="102" swimtime="00:01:58.20" resultid="13160" heatid="14621" lane="4" entrytime="00:02:03.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.80" />
                    <SPLIT distance="50" swimtime="00:00:55.66" />
                    <SPLIT distance="75" swimtime="00:01:27.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="132" swimtime="00:01:28.23" resultid="13161" heatid="14668" lane="2" entrytime="00:01:51.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.53" />
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="75" swimtime="00:01:05.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kassim" lastname="Munshi" birthdate="2007-01-17" gender="M" nation="GBR" license="5701" swrid="4692784" athleteid="13069">
              <RESULTS>
                <RESULT eventid="1117" status="WDR" swimtime="00:00:00.00" resultid="13070" entrytime="00:01:13.74" entrycourse="SCM" />
                <RESULT eventid="1127" status="WDR" swimtime="00:00:00.00" resultid="13071" entrytime="00:01:27.85" entrycourse="SCM" />
                <RESULT eventid="1133" status="WDR" swimtime="00:00:00.00" resultid="13072" entrytime="00:01:04.51" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Muriel" lastname="Zingg" birthdate="2008-03-23" gender="F" nation="SUI" license="32114" swrid="4607541" athleteid="13162">
              <RESULTS>
                <RESULT eventid="1108" points="391" swimtime="00:01:14.65" resultid="13163" heatid="14689" lane="3" entrytime="00:01:17.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.75" />
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="75" swimtime="00:00:54.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="346" swimtime="00:01:18.14" resultid="13164" heatid="14709" lane="2" entrytime="00:01:21.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.22" />
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="75" swimtime="00:00:58.07" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 18:37)" eventid="1124" status="DSQ" swimtime="00:01:23.07" resultid="13165" heatid="14749" lane="1" entrytime="00:01:21.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.56" />
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                    <SPLIT distance="75" swimtime="00:01:00.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="374" swimtime="00:01:09.69" resultid="13166" heatid="14773" lane="2" entrytime="00:01:09.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.50" />
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="75" swimtime="00:00:51.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lionel" lastname="Hofstätter" birthdate="2012-08-07" gender="M" nation="GER" license="32019" swrid="5458190" athleteid="13008">
              <RESULTS>
                <RESULT eventid="1081" points="103" swimtime="00:01:42.93" resultid="13009" heatid="14563" lane="1" entrytime="00:02:01.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.18" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="527 - Wechselbeinschlag während des Schwimmens (Zeit: 12:54)" eventid="1095" status="DSQ" swimtime="00:01:54.57" resultid="13010" heatid="14619" lane="1" entrytime="00:02:06.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.53" />
                    <SPLIT distance="50" swimtime="00:00:53.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="97" swimtime="00:01:37.73" resultid="13011" heatid="14670" lane="3" entrytime="00:01:45.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.11" />
                    <SPLIT distance="50" swimtime="00:00:43.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jayden" lastname="Panzera" birthdate="2011-04-20" gender="M" nation="SUI" license="32022" swrid="5458212" athleteid="13073">
              <RESULTS>
                <RESULT eventid="1071" points="147" swimtime="00:01:30.35" resultid="13074" heatid="14525" lane="1" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.04" />
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                    <SPLIT distance="75" swimtime="00:01:05.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="100" swimtime="00:01:43.80" resultid="13075" heatid="14564" lane="4" entrytime="00:01:57.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.65" />
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                    <SPLIT distance="75" swimtime="00:01:18.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="171" swimtime="00:01:39.60" resultid="13076" heatid="14624" lane="2" entrytime="00:01:50.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.96" />
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                    <SPLIT distance="75" swimtime="00:01:13.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="165" swimtime="00:01:21.80" resultid="13077" heatid="14677" lane="3" entrytime="00:01:26.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.05" />
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="75" swimtime="00:00:59.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celeste" lastname="Kick Bedoya" birthdate="2012-12-30" gender="F" nation="GER" license="21193" swrid="5458197" athleteid="13042">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 9:57)" eventid="1078" status="DSQ" swimtime="00:02:01.56" resultid="13043" heatid="14538" lane="4" entrytime="00:02:37.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.19" />
                    <SPLIT distance="50" swimtime="00:00:56.94" />
                    <SPLIT distance="75" swimtime="00:01:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  2) (Zeit: 12:12)" eventid="1092" status="DSQ" swimtime="00:02:02.24" resultid="13044" heatid="14598" lane="1" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.16" />
                    <SPLIT distance="50" swimtime="00:00:57.86" />
                    <SPLIT distance="75" swimtime="00:01:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="117" swimtime="00:01:42.46" resultid="13045" heatid="14645" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.43" />
                    <SPLIT distance="50" swimtime="00:00:47.58" />
                    <SPLIT distance="75" swimtime="00:01:15.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Rausch" birthdate="2009-07-31" gender="F" nation="SUI" license="5705" swrid="4415949" athleteid="13092">
              <RESULTS>
                <RESULT eventid="1108" points="269" swimtime="00:01:24.52" resultid="13093" heatid="14684" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.55" />
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="75" swimtime="00:00:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="307" swimtime="00:01:21.29" resultid="13094" heatid="14710" lane="2" entrytime="00:01:20.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.95" />
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="75" swimtime="00:01:00.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="323" swimtime="00:01:30.88" resultid="13095" heatid="14745" lane="4" entrytime="00:01:30.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.45" />
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="75" swimtime="00:01:06.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="350" swimtime="00:01:11.28" resultid="13096" heatid="14771" lane="1" entrytime="00:01:12.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.46" />
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="75" swimtime="00:00:53.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lionel" lastname="Jungen" birthdate="2013-05-03" gender="M" nation="SUI" license="5711" swrid="5440823" athleteid="13029">
              <RESULTS>
                <RESULT eventid="1066" points="90" swimtime="00:00:48.39" resultid="13030" heatid="14516" lane="2" entrytime="00:00:51.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="102" swimtime="00:00:47.41" resultid="13031" heatid="14537" lane="2" entrytime="00:00:48.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1090" points="114" swimtime="00:00:51.94" resultid="13032" heatid="14594" lane="2" entrytime="00:00:52.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="133" swimtime="00:00:39.46" resultid="13033" heatid="14641" lane="1" entrytime="00:00:41.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Caddy" birthdate="2008-12-24" gender="F" nation="CZE" license="5663" swrid="5209645" athleteid="12978">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="12979" entrytime="00:01:35.81" entrycourse="SCM" />
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="12980" entrytime="00:01:35.67" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="12981" entrytime="00:01:16.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melanie" lastname="Hutter" birthdate="2009-01-14" gender="F" nation="SUI" license="5733" swrid="4941138" athleteid="13021">
              <RESULTS>
                <RESULT eventid="1114" points="329" swimtime="00:01:19.44" resultid="13022" heatid="14710" lane="4" entrytime="00:01:21.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="75" swimtime="00:01:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="283" swimtime="00:01:34.95" resultid="13023" heatid="14743" lane="3" entrytime="00:01:33.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.69" />
                    <SPLIT distance="50" swimtime="00:00:45.38" />
                    <SPLIT distance="75" swimtime="00:01:10.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="328" swimtime="00:01:12.82" resultid="13024" heatid="14771" lane="4" entrytime="00:01:12.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.63" />
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="75" swimtime="00:00:54.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Shiv" lastname="Thomet" birthdate="2009-02-09" gender="M" nation="SUI" license="32028" swrid="5458167" athleteid="13138">
              <RESULTS>
                <RESULT eventid="1117" points="186" swimtime="00:01:24.57" resultid="13139" heatid="14722" lane="2" entrytime="00:01:23.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="75" swimtime="00:01:03.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="209" swimtime="00:01:33.24" resultid="13140" heatid="14756" lane="3" entrytime="00:01:34.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.72" />
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="75" swimtime="00:01:07.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="231" swimtime="00:01:13.22" resultid="13141" heatid="14786" lane="3" entrytime="00:01:14.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="75" swimtime="00:00:55.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pia" lastname="Salmon" birthdate="2006-09-16" gender="F" nation="GBR" license="5745" swrid="5182839" athleteid="13115">
              <RESULTS>
                <RESULT eventid="1108" points="249" swimtime="00:01:26.73" resultid="13116" heatid="14687" lane="2" entrytime="00:01:25.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.97" />
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                    <SPLIT distance="75" swimtime="00:01:01.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="328" swimtime="00:01:19.53" resultid="13117" heatid="14712" lane="4" entrytime="00:01:17.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.75" />
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Zeit: 18:35)" eventid="1124" status="DSQ" swimtime="00:01:33.05" resultid="13118" heatid="14746" lane="1" entrytime="00:01:28.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.14" />
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                    <SPLIT distance="75" swimtime="00:01:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="336" swimtime="00:01:12.26" resultid="13119" heatid="14773" lane="1" entrytime="00:01:10.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.78" />
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="75" swimtime="00:00:53.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Press" birthdate="2011-07-15" gender="F" nation="SUI" license="5757" swrid="4415959" athleteid="13088">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="13089" entrytime="00:02:02.34" entrycourse="SCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13090" entrytime="00:02:10.37" entrycourse="SCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="13091" entrytime="00:01:49.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matteo" lastname="Baumann" birthdate="2010-05-21" gender="M" nation="SUI" license="5729" swrid="5419460" athleteid="12965">
              <RESULTS>
                <RESULT eventid="1071" points="268" swimtime="00:01:14.06" resultid="12966" heatid="14526" lane="2" entrytime="00:01:12.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.39" />
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="75" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="232" swimtime="00:01:18.55" resultid="12967" heatid="14573" lane="2" entrytime="00:01:17.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.15" />
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="75" swimtime="00:00:58.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="237" swimtime="00:01:29.31" resultid="12968" heatid="14629" lane="3" entrytime="00:01:31.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.25" />
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                    <SPLIT distance="75" swimtime="00:01:06.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="319" swimtime="00:01:05.76" resultid="12969" heatid="14681" lane="2" entrytime="00:01:07.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.78" />
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="75" swimtime="00:00:49.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaja" lastname="Jelinek" birthdate="2012-11-04" gender="F" nation="POL" license="40642" swrid="5508995" athleteid="13025">
              <RESULTS>
                <RESULT eventid="1078" status="DNS" swimtime="00:00:00.00" resultid="13026" heatid="14539" lane="1" entrytime="00:02:12.00" />
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  2) (Zeit: 12:13)" eventid="1092" status="DSQ" swimtime="00:02:02.24" resultid="13027" heatid="14597" lane="1" entrytime="00:02:15.00" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="13028" heatid="14644" lane="3" entrytime="00:02:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Josephine" lastname="Haug" birthdate="2012-04-05" gender="F" nation="SUI" license="32018" swrid="5471570" athleteid="13004">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende 1) (Zeit: 10:00)" eventid="1078" status="DSQ" swimtime="00:01:54.80" resultid="13005" heatid="14540" lane="3" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.83" />
                    <SPLIT distance="50" swimtime="00:00:54.01" />
                    <SPLIT distance="75" swimtime="00:01:24.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="70" swimtime="00:02:30.65" resultid="13006" heatid="14598" lane="4" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.66" />
                    <SPLIT distance="50" swimtime="00:01:08.86" />
                    <SPLIT distance="75" swimtime="00:01:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="107" swimtime="00:01:45.78" resultid="13007" heatid="14645" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.44" />
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                    <SPLIT distance="75" swimtime="00:01:16.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Kaufmann" birthdate="2012-05-09" gender="M" nation="GER" license="21192" swrid="5458196" athleteid="13038">
              <RESULTS>
                <RESULT eventid="1081" points="58" swimtime="00:02:04.18" resultid="13039" heatid="14561" lane="4" entrytime="00:02:06.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.96" />
                    <SPLIT distance="50" swimtime="00:00:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="95" swimtime="00:02:01.15" resultid="13040" heatid="14619" lane="4" entrytime="00:02:07.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.48" />
                    <SPLIT distance="50" swimtime="00:00:56.07" />
                    <SPLIT distance="75" swimtime="00:01:28.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="75" swimtime="00:01:46.15" resultid="13041" heatid="14670" lane="4" entrytime="00:01:48.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.15" />
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                    <SPLIT distance="75" swimtime="00:01:17.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulina" lastname="Roth" birthdate="2006-11-16" gender="F" nation="SUI" license="5744" swrid="4415954" athleteid="13108">
              <RESULTS>
                <RESULT eventid="1124" points="253" swimtime="00:01:38.47" resultid="13109" heatid="14741" lane="3" entrytime="00:01:39.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.87" />
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                    <SPLIT distance="75" swimtime="00:01:12.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="287" swimtime="00:01:16.18" resultid="13110" heatid="14769" lane="1" entrytime="00:01:16.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.47" />
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="75" swimtime="00:00:57.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yeholy" lastname="Schwartz" birthdate="2008-08-22" gender="F" nation="SUI" license="42480" swrid="5309714" athleteid="13125">
              <RESULTS>
                <RESULT eventid="1114" points="179" swimtime="00:01:37.26" resultid="13126" heatid="14704" lane="2" entrytime="00:01:35.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:12.60" />
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="194" swimtime="00:01:47.71" resultid="13127" heatid="14739" lane="2" entrytime="00:01:48.87">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.97" />
                    <SPLIT distance="50" swimtime="00:00:50.04" />
                    <SPLIT distance="75" swimtime="00:01:18.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="161" swimtime="00:01:32.19" resultid="13128" heatid="14765" lane="2" entrytime="00:01:28.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.08" />
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                    <SPLIT distance="75" swimtime="00:01:08.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatrice" lastname="Cussigh" birthdate="2007-04-28" gender="F" nation="SUI" license="5669" swrid="4040977" athleteid="12987">
              <RESULTS>
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="12988" heatid="14691" lane="2" entrytime="00:01:11.25" entrycourse="SCM" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="12989" heatid="14711" lane="3" entrytime="00:01:18.23" entrycourse="SCM" />
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="12990" heatid="14780" lane="4" entrytime="00:01:02.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henri" lastname="Siegmann" birthdate="2012-03-03" gender="M" nation="GER" athleteid="13129">
              <RESULTS>
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene (Zeit: 12:43)" eventid="1095" status="DSQ" swimtime="00:02:22.01" resultid="13130" heatid="14615" lane="1" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.89" />
                    <SPLIT distance="50" swimtime="00:01:06.97" />
                    <SPLIT distance="75" swimtime="00:01:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="58" swimtime="00:01:55.55" resultid="13131" heatid="14665" lane="2" entrytime="00:02:12.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.27" />
                    <SPLIT distance="50" swimtime="00:00:55.68" />
                    <SPLIT distance="75" swimtime="00:01:27.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="51" swimtime="00:02:09.87" resultid="13132" heatid="14559" lane="1" entrytime="00:02:25.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.37" />
                    <SPLIT distance="50" swimtime="00:01:02.15" />
                    <SPLIT distance="75" swimtime="00:01:36.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Aufdereggen" birthdate="2010-07-26" gender="F" nation="SUI" license="5679" swrid="5351140" athleteid="12961">
              <RESULTS>
                <RESULT eventid="1078" points="181" swimtime="00:01:36.91" resultid="12962" heatid="14550" lane="1" entrytime="00:01:36.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.14" />
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="75" swimtime="00:01:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="231" swimtime="00:01:41.49" resultid="12963" heatid="14606" lane="4" entrytime="00:01:43.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.69" />
                    <SPLIT distance="50" swimtime="00:00:47.12" />
                    <SPLIT distance="75" swimtime="00:01:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="234" swimtime="00:01:21.52" resultid="12964" heatid="14658" lane="1" entrytime="00:01:21.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.26" />
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                    <SPLIT distance="75" swimtime="00:01:00.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tamara" lastname="Braschler" birthdate="2012-01-06" gender="F" nation="SUI" license="5760" swrid="5440818" athleteid="12974">
              <RESULTS>
                <RESULT eventid="1078" points="119" swimtime="00:01:51.47" resultid="12975" heatid="14542" lane="2" entrytime="00:01:55.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.72" />
                    <SPLIT distance="50" swimtime="00:00:54.02" />
                    <SPLIT distance="75" swimtime="00:01:24.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="181" swimtime="00:01:50.20" resultid="12976" heatid="14602" lane="4" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.42" />
                    <SPLIT distance="50" swimtime="00:00:51.95" />
                    <SPLIT distance="75" swimtime="00:01:21.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="125" swimtime="00:01:40.38" resultid="12977" heatid="14650" lane="2" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.98" />
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="75" swimtime="00:01:15.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Collin" lastname="Schmidlin" birthdate="2001-03-21" gender="M" nation="SUI" license="5672" swrid="4777365" athleteid="13120" />
            <ATHLETE firstname="Aksel" lastname="Just" birthdate="2012-04-03" gender="M" nation="DEN" license="38116" swrid="5489036" athleteid="13034">
              <RESULTS>
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="13035" entrytime="00:01:55.00" />
                <RESULT eventid="1095" status="WDR" swimtime="00:00:00.00" resultid="13036" entrytime="00:02:10.94" entrycourse="LCM" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="13037" entrytime="00:01:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Finn" lastname="Rieger" birthdate="2007-04-25" gender="M" nation="GER" license="5686" swrid="5340078" athleteid="13100">
              <RESULTS>
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="13101" entrytime="00:01:15.09" entrycourse="SCM" />
                <RESULT eventid="1117" status="WDR" swimtime="00:00:00.00" resultid="13102" entrytime="00:01:22.05" entrycourse="SCM" />
                <RESULT eventid="1133" status="WDR" swimtime="00:00:00.00" resultid="13103" entrytime="00:01:04.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estrid" lastname="Wittner" birthdate="2009-11-27" gender="F" nation="SWE" license="40207" swrid="5503642" athleteid="13150">
              <RESULTS>
                <RESULT eventid="1114" points="140" swimtime="00:01:45.55" resultid="13151" heatid="14703" lane="2" entrytime="00:01:45.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.44" />
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="220" swimtime="00:01:43.24" resultid="13152" heatid="14739" lane="1" entrytime="00:01:54.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.50" />
                    <SPLIT distance="50" swimtime="00:00:48.22" />
                    <SPLIT distance="75" swimtime="00:01:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="135" swimtime="00:01:37.83" resultid="13153" heatid="14765" lane="1" entrytime="00:01:42.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.43" />
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                    <SPLIT distance="75" swimtime="00:01:12.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Woods" birthdate="2012-09-06" gender="F" nation="AUT" license="40637" swrid="5509030" athleteid="13154">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende 1) (Zeit: 9:57)" eventid="1078" status="DSQ" swimtime="00:02:04.27" resultid="13155" heatid="14538" lane="3" entrytime="00:02:26.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.21" />
                    <SPLIT distance="50" swimtime="00:01:00.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="67" swimtime="00:02:32.80" resultid="13156" heatid="14595" lane="3" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.33" />
                    <SPLIT distance="50" swimtime="00:01:10.54" />
                    <SPLIT distance="75" swimtime="00:01:52.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="98" swimtime="00:01:48.71" resultid="13157" heatid="14643" lane="3" entrytime="00:02:19.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.96" />
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                    <SPLIT distance="75" swimtime="00:01:18.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luise" lastname="Robrahn" birthdate="2012-12-13" gender="F" nation="GER" license="21197" swrid="5458215" athleteid="13104">
              <RESULTS>
                <RESULT eventid="1078" points="82" swimtime="00:02:06.11" resultid="13105" heatid="14541" lane="1" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.67" />
                    <SPLIT distance="50" swimtime="00:00:59.27" />
                    <SPLIT distance="75" swimtime="00:01:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="136" swimtime="00:02:01.24" resultid="13106" heatid="14600" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.52" />
                    <SPLIT distance="50" swimtime="00:00:56.41" />
                    <SPLIT distance="75" swimtime="00:01:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="102" swimtime="00:01:47.51" resultid="13107" heatid="14646" lane="1" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.99" />
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="75" swimtime="00:01:19.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anouk" lastname="Schumacher" birthdate="2008-02-01" gender="F" nation="SUI" license="5665" swrid="5419463" athleteid="13121">
              <RESULTS>
                <RESULT eventid="1114" points="141" swimtime="00:01:45.34" resultid="13122" heatid="14704" lane="3" entrytime="00:01:43.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="169" swimtime="00:01:52.77" resultid="13123" heatid="14739" lane="3" entrytime="00:01:49.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.61" />
                    <SPLIT distance="50" swimtime="00:00:52.86" />
                    <SPLIT distance="75" swimtime="00:01:22.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="197" swimtime="00:01:26.33" resultid="13124" heatid="14766" lane="1" entrytime="00:01:28.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.51" />
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="75" swimtime="00:01:05.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luca" lastname="Rusu" birthdate="2012-05-12" gender="M" nation="SUI" license="32025" swrid="5458216" athleteid="13111">
              <RESULTS>
                <RESULT eventid="1081" points="51" swimtime="00:02:09.94" resultid="13112" heatid="14559" lane="3" entrytime="00:02:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.77" />
                    <SPLIT distance="50" swimtime="00:01:01.95" />
                    <SPLIT distance="75" swimtime="00:01:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="77" swimtime="00:02:09.97" resultid="13113" heatid="14616" lane="1" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.13" />
                    <SPLIT distance="50" swimtime="00:01:02.09" />
                    <SPLIT distance="75" swimtime="00:01:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="43" swimtime="00:02:08.13" resultid="13114" heatid="14667" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.14" />
                    <SPLIT distance="50" swimtime="00:00:58.44" />
                    <SPLIT distance="75" swimtime="00:01:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Malcolm" lastname="Mensah" birthdate="2006-02-23" gender="M" nation="SUI" license="5718" swrid="5092502" athleteid="13066">
              <RESULTS>
                <RESULT eventid="1127" points="283" swimtime="00:01:24.25" resultid="13067" heatid="14760" lane="4" entrytime="00:01:22.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.88" />
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="75" swimtime="00:01:01.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="322" swimtime="00:01:05.50" resultid="13068" heatid="14790" lane="2" entrytime="00:01:04.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.69" />
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="75" swimtime="00:00:49.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elena" lastname="Meili" birthdate="2010-12-25" gender="F" nation="SUI" license="5676" swrid="5351149" athleteid="13054">
              <RESULTS>
                <RESULT eventid="1078" points="145" swimtime="00:01:44.32" resultid="13055" heatid="14546" lane="2" entrytime="00:01:44.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.85" />
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="209" swimtime="00:01:44.93" resultid="13056" heatid="14604" lane="3" entrytime="00:01:48.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.61" />
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                    <SPLIT distance="75" swimtime="00:01:16.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="181" swimtime="00:01:28.83" resultid="13057" heatid="14651" lane="2" entrytime="00:01:31.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:04.69" />
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Louan" lastname="Brand" birthdate="2009-01-06" gender="M" nation="SUI" license="5713" swrid="5419461" athleteid="12970">
              <RESULTS>
                <RESULT eventid="1117" points="134" swimtime="00:01:34.37" resultid="12971" heatid="14722" lane="4" entrytime="00:01:25.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.80" />
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="75" swimtime="00:01:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="145" swimtime="00:01:45.15" resultid="12972" heatid="14754" lane="3" entrytime="00:01:45.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.06" />
                    <SPLIT distance="50" swimtime="00:00:49.62" />
                    <SPLIT distance="75" swimtime="00:01:17.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="218" swimtime="00:01:14.66" resultid="12973" heatid="14786" lane="1" entrytime="00:01:15.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="75" swimtime="00:00:55.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Wienecke" birthdate="2011-07-05" gender="F" nation="GER" license="5743" swrid="5382441" athleteid="13146">
              <RESULTS>
                <RESULT eventid="1078" points="145" swimtime="00:01:44.28" resultid="13147" heatid="14543" lane="1" entrytime="00:01:51.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.08" />
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="75" swimtime="00:01:19.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="195" swimtime="00:01:47.47" resultid="13148" heatid="14599" lane="4" entrytime="00:02:07.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.38" />
                    <SPLIT distance="50" swimtime="00:00:49.85" />
                    <SPLIT distance="75" swimtime="00:01:18.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="193" swimtime="00:01:26.88" resultid="13149" heatid="14653" lane="1" entrytime="00:01:27.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="75" swimtime="00:01:03.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer 2) (Zeit: 11:38)" eventid="1086" status="DSQ" swimtime="00:02:24.90" resultid="13167" heatid="14818" lane="1" entrytime="00:02:16.93">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.07" />
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                    <SPLIT distance="75" swimtime="00:00:58.00" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="125" swimtime="00:01:36.02" />
                    <SPLIT distance="150" swimtime="00:01:55.65" />
                    <SPLIT distance="175" swimtime="00:02:09.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13029" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="13158" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="13073" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="12965" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="300" swimtime="00:02:15.02" resultid="13168" heatid="14735" lane="2" entrytime="00:02:07.64">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.60" />
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="75" swimtime="00:00:52.53" />
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                    <SPLIT distance="125" swimtime="00:01:26.79" />
                    <SPLIT distance="150" swimtime="00:01:43.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12996" number="1" />
                    <RELAYPOSITION athleteid="13066" number="2" />
                    <RELAYPOSITION athleteid="13120" number="3" />
                    <RELAYPOSITION athleteid="13097" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1086" points="87" swimtime="00:03:04.13" resultid="13169" heatid="14583" lane="1" entrytime="00:02:39.28">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.21" />
                    <SPLIT distance="50" swimtime="00:00:57.37" />
                    <SPLIT distance="75" swimtime="00:01:17.16" />
                    <SPLIT distance="100" swimtime="00:01:39.75" />
                    <SPLIT distance="125" swimtime="00:01:59.70" />
                    <SPLIT distance="150" swimtime="00:02:23.89" />
                    <SPLIT distance="175" swimtime="00:02:42.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13111" number="1" />
                    <RELAYPOSITION athleteid="13008" number="2" />
                    <RELAYPOSITION athleteid="13038" number="3" />
                    <RELAYPOSITION athleteid="13050" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1122" status="WDR" swimtime="00:00:00.00" resultid="13170" entrytime="00:02:20.91">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13097" number="1" />
                    <RELAYPOSITION athleteid="13069" number="2" />
                    <RELAYPOSITION athleteid="13100" number="3" />
                    <RELAYPOSITION athleteid="13058" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="246" swimtime="00:02:27.43" resultid="13171" heatid="14580" lane="3" entrytime="00:02:28.26">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.67" />
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="75" swimtime="00:00:54.57" />
                    <SPLIT distance="100" swimtime="00:01:13.66" />
                    <SPLIT distance="125" swimtime="00:01:30.84" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                    <SPLIT distance="175" swimtime="00:02:07.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13012" number="1" />
                    <RELAYPOSITION athleteid="13016" number="2" />
                    <RELAYPOSITION athleteid="13054" number="3" />
                    <RELAYPOSITION athleteid="13078" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="391" swimtime="00:02:19.92" resultid="13172" heatid="14732" lane="2" entrytime="00:02:12.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="75" swimtime="00:00:54.92" />
                    <SPLIT distance="100" swimtime="00:01:15.93" />
                    <SPLIT distance="125" swimtime="00:01:31.85" />
                    <SPLIT distance="150" swimtime="00:01:51.86" />
                    <SPLIT distance="175" swimtime="00:02:05.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13115" number="1" />
                    <RELAYPOSITION athleteid="13162" number="2" />
                    <RELAYPOSITION athleteid="13092" number="3" />
                    <RELAYPOSITION athleteid="13083" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer 4) (Zeit: 11:16)" eventid="1084" status="DSQ" swimtime="00:02:37.97" resultid="13173" heatid="14579" lane="3" entrytime="00:02:38.17">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.79" />
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                    <SPLIT distance="75" swimtime="00:00:56.97" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="125" swimtime="00:01:39.02" />
                    <SPLIT distance="150" swimtime="00:02:02.32" />
                    <SPLIT distance="175" swimtime="00:02:18.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13146" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="12974" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="12956" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="12961" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1120" points="309" swimtime="00:02:31.43" resultid="13174" heatid="14731" lane="3" entrytime="00:02:35.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.99" />
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                    <SPLIT distance="75" swimtime="00:00:56.58" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="125" swimtime="00:01:37.38" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                    <SPLIT distance="175" swimtime="00:02:14.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13021" number="1" />
                    <RELAYPOSITION athleteid="13000" number="2" />
                    <RELAYPOSITION athleteid="13142" number="3" />
                    <RELAYPOSITION athleteid="13108" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1084" points="125" swimtime="00:03:04.91" resultid="13175" heatid="14578" lane="4" entrytime="00:02:54.76">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.78" />
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="75" swimtime="00:01:06.39" />
                    <SPLIT distance="100" swimtime="00:01:32.32" />
                    <SPLIT distance="125" swimtime="00:01:53.50" />
                    <SPLIT distance="150" swimtime="00:02:20.51" />
                    <SPLIT distance="175" swimtime="00:02:41.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13042" number="1" />
                    <RELAYPOSITION athleteid="13154" number="2" />
                    <RELAYPOSITION athleteid="13104" number="3" />
                    <RELAYPOSITION athleteid="13004" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="FTAL" nation="SUI" region="RZW" clubid="13393" swrid="65685" name="Schwimmclub Fricktal">
          <ATHLETES>
            <ATHLETE firstname="Helena" lastname="Krzeminska" birthdate="2011-04-28" gender="F" nation="POL" license="35580" swrid="4856046" athleteid="13914">
              <RESULTS>
                <RESULT eventid="1078" points="124" swimtime="00:01:49.93" resultid="13915" heatid="14542" lane="3" entrytime="00:01:56.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:01:21.38" />
                    <SPLIT distance="50" swimtime="00:00:52.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="109" swimtime="00:02:10.38" resultid="13916" heatid="14596" lane="4" entrytime="00:02:24.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.96" />
                    <SPLIT distance="50" swimtime="00:01:00.78" />
                    <SPLIT distance="75" swimtime="00:01:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="138" swimtime="00:01:37.03" resultid="13917" heatid="14646" lane="2" entrytime="00:01:47.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.24" />
                    <SPLIT distance="50" swimtime="00:00:46.31" />
                    <SPLIT distance="75" swimtime="00:01:13.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Nikolic" birthdate="2012-01-01" gender="F" nation="SUI" license="34949" swrid="4856303" athleteid="13927">
              <RESULTS>
                <RESULT eventid="1078" points="156" swimtime="00:01:41.82" resultid="13928" heatid="14545" lane="1" entrytime="00:01:46.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.71" />
                    <SPLIT distance="50" swimtime="00:00:50.94" />
                    <SPLIT distance="75" swimtime="00:01:16.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="135" swimtime="00:02:01.45" resultid="13929" heatid="14599" lane="2" entrytime="00:02:05.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.89" />
                    <SPLIT distance="50" swimtime="00:00:56.99" />
                    <SPLIT distance="75" swimtime="00:01:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="123" swimtime="00:01:40.84" resultid="13930" heatid="14650" lane="3" entrytime="00:01:37.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.27" />
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                    <SPLIT distance="75" swimtime="00:01:17.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Eiselt" birthdate="2014-11-17" gender="F" nation="SUI" license="40215" swrid="5523263" athleteid="13869">
              <RESULTS>
                <RESULT eventid="1074" points="81" swimtime="00:00:58.96" resultid="13870" heatid="14530" lane="4" entrytime="00:01:02.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:28.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="95" swimtime="00:01:02.48" resultid="13871" heatid="14587" lane="2" entrytime="00:01:05.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="90" swimtime="00:00:51.12" resultid="13872" heatid="14634" lane="4" entrytime="00:00:58.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Debora" lastname="Mettler" birthdate="2011-05-06" gender="F" nation="SUI" license="7602" swrid="5365450" athleteid="13918">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="13919" entrytime="00:01:54.54" entrycourse="SCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13920" entrytime="00:02:01.39" entrycourse="LCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="13921" entrytime="00:01:29.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mona" lastname="Wetli" birthdate="2013-04-06" gender="F" nation="SUI" license="40212" swrid="5523273" athleteid="13965">
              <RESULTS>
                <RESULT eventid="1074" points="81" swimtime="00:00:58.97" resultid="13966" heatid="14529" lane="4" entrytime="00:01:07.28" entrycourse="SCM" />
                <RESULT eventid="1088" points="70" swimtime="00:01:09.04" resultid="13967" heatid="14585" lane="1" entrytime="00:01:18.35" entrycourse="LCM" />
                <RESULT eventid="1098" points="96" swimtime="00:00:50.05" resultid="13968" heatid="14633" lane="4" entrytime="00:01:02.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raya" lastname="Benz" birthdate="2014-03-05" gender="F" nation="SUI" license="34938" swrid="4854385" athleteid="13851">
              <RESULTS>
                <RESULT eventid="1074" points="81" swimtime="00:00:59.14" resultid="13852" heatid="14531" lane="4" entrytime="00:00:59.98" entrycourse="SCM" />
                <RESULT eventid="1088" points="46" swimtime="00:01:19.21" resultid="13853" heatid="14584" lane="3" entrytime="00:01:21.87" entrycourse="SCM" />
                <RESULT eventid="1098" points="42" swimtime="00:01:05.71" resultid="13854" heatid="14632" lane="2" entrytime="00:01:03.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Kovac" birthdate="2012-08-02" gender="M" nation="SUI" license="34936" swrid="4855992" athleteid="13908">
              <RESULTS>
                <RESULT eventid="1081" points="69" swimtime="00:01:57.72" resultid="13909" heatid="14559" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.40" />
                    <SPLIT distance="50" swimtime="00:00:58.70" />
                    <SPLIT distance="75" swimtime="00:01:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="42" swimtime="00:02:08.42" resultid="13910" heatid="14666" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.12" />
                    <SPLIT distance="50" swimtime="00:00:58.70" />
                    <SPLIT distance="75" swimtime="00:01:33.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julius" lastname="Ilten" birthdate="2004-01-23" gender="M" nation="GER" license="7616" swrid="5105411" athleteid="13903">
              <RESULTS>
                <RESULT eventid="1111" points="359" swimtime="00:01:07.21" resultid="13904" heatid="14698" lane="2" entrytime="00:01:08.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.46" />
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                    <SPLIT distance="75" swimtime="00:00:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="390" swimtime="00:01:06.10" resultid="13905" heatid="14728" lane="1" entrytime="00:01:05.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.54" />
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="75" swimtime="00:00:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="397" swimtime="00:01:15.26" resultid="13906" heatid="14762" lane="3" entrytime="00:01:11.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.31" />
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="75" swimtime="00:00:55.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="455" swimtime="00:00:58.41" resultid="13907" heatid="14795" lane="2" entrytime="00:00:56.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.21" />
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="75" swimtime="00:00:43.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Gisler" birthdate="2006-07-29" gender="F" nation="SUI" license="7629" swrid="5278961" athleteid="13891">
              <RESULTS>
                <RESULT eventid="1114" points="409" swimtime="00:01:13.92" resultid="13892" heatid="14712" lane="1" entrytime="00:01:17.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.04" />
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="75" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="333" swimtime="00:01:29.89" resultid="13893" heatid="14746" lane="3" entrytime="00:01:28.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.85" />
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="75" swimtime="00:01:05.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="486" swimtime="00:01:03.87" resultid="13894" heatid="14777" lane="4" entrytime="00:01:05.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.22" />
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                    <SPLIT distance="75" swimtime="00:00:46.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lewis" lastname="Rippstein" birthdate="2006-01-02" gender="M" nation="SUI" license="7620" swrid="5053849" athleteid="13931">
              <RESULTS>
                <RESULT eventid="1111" points="445" swimtime="00:01:02.58" resultid="13932" heatid="14700" lane="1" entrytime="00:01:03.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.99" />
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                    <SPLIT distance="75" swimtime="00:00:45.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="356" swimtime="00:01:08.16" resultid="13933" heatid="14727" lane="3" entrytime="00:01:08.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.70" />
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="75" swimtime="00:00:50.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="331" swimtime="00:01:19.97" resultid="13934" heatid="14761" lane="1" entrytime="00:01:17.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.58" />
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                    <SPLIT distance="75" swimtime="00:00:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="499" swimtime="00:00:56.65" resultid="13935" heatid="14795" lane="1" entrytime="00:00:56.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:12.60" />
                    <SPLIT distance="50" swimtime="00:00:26.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Linda" lastname="Egger" birthdate="2007-08-15" gender="F" nation="SUI" license="7623" swrid="5157248" athleteid="13864">
              <RESULTS>
                <RESULT eventid="1108" points="371" swimtime="00:01:15.99" resultid="13865" heatid="14689" lane="1" entrytime="00:01:17.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.30" />
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="75" swimtime="00:00:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="475" swimtime="00:01:10.33" resultid="13866" heatid="14715" lane="2" entrytime="00:01:09.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.51" />
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="75" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="386" swimtime="00:01:25.61" resultid="13867" heatid="14745" lane="2" entrytime="00:01:29.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="75" swimtime="00:01:02.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="526" swimtime="00:01:02.24" resultid="13868" heatid="14780" lane="2" entrytime="00:01:01.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.25" />
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="75" swimtime="00:00:46.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6685" points="481" swimtime="00:00:32.66" resultid="14847" heatid="14801" lane="4" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roman" lastname="Strashnov" birthdate="2011-07-01" gender="M" nation="GER" athleteid="13944">
              <RESULTS>
                <RESULT eventid="1081" points="63" swimtime="00:02:00.86" resultid="13945" heatid="14562" lane="1" entrytime="00:02:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                    <SPLIT distance="75" swimtime="00:01:27.95" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="999 - , 113 - Rennen nicht beendet" eventid="1105" status="DSQ" swimtime="00:02:22.23" resultid="13946" heatid="14668" lane="4" entrytime="00:01:58.01">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.24" />
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="75" swimtime="00:01:20.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Sutter" birthdate="2007-04-16" gender="F" nation="SUI" license="7596" swrid="5157250" athleteid="13947">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="13948" entrytime="00:01:24.78" entrycourse="SCM" />
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="13949" entrytime="00:01:22.75" entrycourse="SCM" />
                <RESULT eventid="1124" status="WDR" swimtime="00:00:00.00" resultid="13950" entrytime="00:01:33.71" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="13951" entrytime="00:01:07.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lukas" lastname="Berzins" birthdate="2013-02-25" gender="M" nation="SUI" license="40216" swrid="5540953" athleteid="13855">
              <RESULTS>
                <RESULT eventid="1076" status="WDR" swimtime="00:00:00.00" resultid="13856" entrytime="00:01:04.00" />
                <RESULT eventid="1090" status="WDR" swimtime="00:00:00.00" resultid="13857" entrytime="00:01:10.09" entrycourse="SCM" />
                <RESULT eventid="1100" status="WDR" swimtime="00:00:00.00" resultid="13858" entrytime="00:00:56.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lamar" lastname="Horani" birthdate="2013-07-09" gender="F" nation="SUI" license="40214" swrid="5523264" athleteid="13899">
              <RESULTS>
                <RESULT eventid="1064" points="55" swimtime="00:01:04.06" resultid="13900" heatid="14513" lane="1" entrytime="00:01:01.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.53" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...) (Zeit: 9:17)" eventid="1074" status="DSQ" swimtime="00:00:54.67" resultid="13901" heatid="14531" lane="3" entrytime="00:00:59.90">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="127" swimtime="00:00:45.53" resultid="13902" heatid="14636" lane="3" entrytime="00:00:47.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konstantin" lastname="Stikhin" birthdate="2010-12-14" gender="M" nation="SUI" license="35173" swrid="4856382" athleteid="13941">
              <RESULTS>
                <RESULT eventid="1081" points="50" swimtime="00:02:10.74" resultid="13942" heatid="14560" lane="3" entrytime="00:02:08.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.65" />
                    <SPLIT distance="50" swimtime="00:01:02.41" />
                    <SPLIT distance="75" swimtime="00:01:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando (Zeit: 14:25)" eventid="1105" status="DSQ" swimtime="00:02:05.99" resultid="13943" heatid="14666" lane="1" entrytime="00:02:09.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.76" />
                    <SPLIT distance="50" swimtime="00:00:55.69" />
                    <SPLIT distance="75" swimtime="00:01:33.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nela" lastname="Hanak" birthdate="2012-04-12" gender="F" nation="SUI" license="7630" swrid="5382477" athleteid="13895">
              <RESULTS>
                <RESULT eventid="1078" points="155" swimtime="00:01:42.11" resultid="13896" heatid="14548" lane="2" entrytime="00:01:40.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="192" swimtime="00:01:47.98" resultid="13897" heatid="14604" lane="1" entrytime="00:01:49.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:22.43" />
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                    <SPLIT distance="75" swimtime="00:01:18.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="142" swimtime="00:01:36.12" resultid="13898" heatid="14649" lane="1" entrytime="00:01:39.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.54" />
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jolina" lastname="Wächter" birthdate="2004-07-10" gender="F" nation="SUI" license="7612" swrid="4879743" athleteid="13960">
              <RESULTS>
                <RESULT eventid="1108" points="323" swimtime="00:01:19.56" resultid="13961" heatid="14690" lane="2" entrytime="00:01:14.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.95" />
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="75" swimtime="00:00:57.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="322" swimtime="00:01:20.03" resultid="13962" heatid="14713" lane="4" entrytime="00:01:16.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="271" swimtime="00:01:36.36" resultid="13963" heatid="14743" lane="1" entrytime="00:01:33.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.41" />
                    <SPLIT distance="50" swimtime="00:00:44.89" />
                    <SPLIT distance="75" swimtime="00:01:10.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="357" swimtime="00:01:10.82" resultid="13964" heatid="14775" lane="3" entrytime="00:01:07.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.76" />
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="75" swimtime="00:00:52.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amélie" lastname="Friesewinkel" birthdate="2011-02-04" gender="F" nation="SUI" license="19944" swrid="5440437" athleteid="13873">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="13874" entrytime="00:01:54.49" entrycourse="LCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13875" entrytime="00:01:54.46" entrycourse="LCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="13876" entrytime="00:01:29.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrin" lastname="Gallert" birthdate="2009-08-07" gender="M" nation="SUI" license="7590" swrid="4918220" athleteid="13877">
              <RESULTS>
                <RESULT eventid="1111" points="124" swimtime="00:01:35.67" resultid="13878" heatid="14695" lane="2" entrytime="00:01:34.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.78" />
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                    <SPLIT distance="75" swimtime="00:01:07.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="182" swimtime="00:01:25.19" resultid="13879" heatid="14720" lane="1" entrytime="00:01:37.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.00" />
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="75" swimtime="00:01:03.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="199" swimtime="00:01:34.73" resultid="13880" heatid="14755" lane="1" entrytime="00:01:37.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.78" />
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                    <SPLIT distance="75" swimtime="00:01:11.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="224" swimtime="00:01:13.89" resultid="13881" heatid="14785" lane="2" entrytime="00:01:15.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.27" />
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="75" swimtime="00:00:54.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noa" lastname="Sutter" birthdate="2010-08-05" gender="M" nation="SUI" license="7635" swrid="5326523" athleteid="13952">
              <RESULTS>
                <RESULT eventid="1081" points="76" swimtime="00:01:53.78" resultid="13953" heatid="14566" lane="4" entrytime="00:01:49.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.40" />
                    <SPLIT distance="50" swimtime="00:00:53.61" />
                    <SPLIT distance="75" swimtime="00:01:23.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="125" swimtime="00:01:50.62" resultid="13954" heatid="14625" lane="3" entrytime="00:01:49.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.03" />
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                    <SPLIT distance="75" swimtime="00:01:20.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="98" swimtime="00:01:37.30" resultid="13955" heatid="14671" lane="2" entrytime="00:01:39.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.60" />
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="75" swimtime="00:01:12.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Traver" lastname="Dinten" birthdate="2004-09-28" gender="M" nation="SUI" license="34965" swrid="4830859" athleteid="13859">
              <RESULTS>
                <RESULT eventid="1111" points="414" swimtime="00:01:04.06" resultid="13860" heatid="14699" lane="3" entrytime="00:01:05.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.20" />
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                    <SPLIT distance="75" swimtime="00:00:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="394" swimtime="00:01:05.88" resultid="13861" heatid="14725" lane="1" entrytime="00:01:12.80">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.53" />
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                    <SPLIT distance="75" swimtime="00:00:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="394" swimtime="00:01:15.45" resultid="13862" heatid="14760" lane="2" entrytime="00:01:18.02">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.22" />
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="75" swimtime="00:00:55.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="469" swimtime="00:00:57.82" resultid="13863" heatid="14792" lane="3" entrytime="00:01:00.92">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.25" />
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                    <SPLIT distance="75" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliette" lastname="Siegfried" birthdate="2008-04-11" gender="F" nation="SUI" license="7615" swrid="5157249" athleteid="13936">
              <RESULTS>
                <RESULT eventid="1108" points="357" swimtime="00:01:16.98" resultid="13937" heatid="14690" lane="3" entrytime="00:01:14.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.28" />
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="75" swimtime="00:00:54.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="396" swimtime="00:01:14.71" resultid="13938" heatid="14714" lane="1" entrytime="00:01:13.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.16" />
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="75" swimtime="00:00:55.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="431" swimtime="00:01:22.54" resultid="13939" heatid="14749" lane="4" entrytime="00:01:21.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.44" />
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="75" swimtime="00:01:00.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="432" swimtime="00:01:06.43" resultid="13940" heatid="14777" lane="3" entrytime="00:01:05.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.36" />
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="75" swimtime="00:00:48.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric Keizo" lastname="Tomita" birthdate="2012-05-01" gender="M" nation="GER" license="19946" swrid="5440451" athleteid="13956">
              <RESULTS>
                <RESULT eventid="1081" points="70" swimtime="00:01:56.99" resultid="13957" heatid="14562" lane="3" entrytime="00:02:01.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:27.10" />
                    <SPLIT distance="50" swimtime="00:00:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="82" swimtime="00:02:06.96" resultid="13958" heatid="14620" lane="4" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.96" />
                    <SPLIT distance="50" swimtime="00:00:58.50" />
                    <SPLIT distance="75" swimtime="00:01:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="100" swimtime="00:01:36.62" resultid="13959" heatid="14671" lane="4" entrytime="00:01:40.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.64" />
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="75" swimtime="00:01:13.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elina" lastname="Gallert" birthdate="2007-05-12" gender="F" nation="SUI" license="7603" swrid="5105410" athleteid="13882">
              <RESULTS>
                <RESULT eventid="1108" points="268" swimtime="00:01:24.63" resultid="13883" heatid="14688" lane="3" entrytime="00:01:22.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.25" />
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="75" swimtime="00:01:00.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="330" swimtime="00:01:19.38" resultid="13884" heatid="14707" lane="3" entrytime="00:01:26.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.56" />
                    <SPLIT distance="50" swimtime="00:00:38.30" />
                    <SPLIT distance="75" swimtime="00:00:58.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="324" swimtime="00:01:30.79" resultid="13885" heatid="14745" lane="3" entrytime="00:01:29.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.70" />
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="75" swimtime="00:01:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="355" swimtime="00:01:10.92" resultid="13886" heatid="14774" lane="4" entrytime="00:01:09.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.61" />
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="75" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilia" lastname="Krzeminska" birthdate="2014-10-04" gender="F" nation="POL" license="36945" swrid="5481974" athleteid="13911">
              <RESULTS>
                <RESULT eventid="1074" points="58" swimtime="00:01:05.79" resultid="13912" heatid="14528" lane="3" entrytime="00:01:10.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="47" swimtime="00:01:03.46" resultid="13913" heatid="14631" lane="2" entrytime="00:01:13.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlon" lastname="Mühlebach" birthdate="2006-02-09" gender="M" nation="SUI" license="42211" swrid="5053834" athleteid="13922">
              <RESULTS>
                <RESULT eventid="1111" points="331" swimtime="00:01:09.01" resultid="13923" heatid="14698" lane="1" entrytime="00:01:10.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.34" />
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="75" swimtime="00:00:49.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="321" swimtime="00:01:10.56" resultid="13924" heatid="14725" lane="2" entrytime="00:01:12.24">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.16" />
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="75" swimtime="00:00:52.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="461" swimtime="00:01:11.62" resultid="13925" heatid="14762" lane="4" entrytime="00:01:12.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.42" />
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="75" swimtime="00:00:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="416" swimtime="00:01:00.18" resultid="13926" heatid="14794" lane="4" entrytime="00:00:59.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.54" />
                    <SPLIT distance="50" swimtime="00:00:28.37" />
                    <SPLIT distance="75" swimtime="00:00:44.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arik" lastname="Benz" birthdate="2012-06-05" gender="M" nation="SUI" license="7594" swrid="5425621" athleteid="13847">
              <RESULTS>
                <RESULT eventid="1071" status="WDR" swimtime="00:00:00.00" resultid="13848" entrytime="00:01:35.57" entrycourse="SCM" />
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="13849" entrytime="00:01:48.00" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="13850" entrytime="00:01:25.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norina" lastname="Gallert" birthdate="2011-12-11" gender="F" nation="SUI" license="7636" swrid="5353511" athleteid="13887">
              <RESULTS>
                <RESULT eventid="1078" status="WDR" swimtime="00:00:00.00" resultid="13888" entrytime="00:02:09.70" entrycourse="SCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13889" entrytime="00:01:59.78" entrycourse="SCM" />
                <RESULT eventid="1102" status="WDR" swimtime="00:00:00.00" resultid="13890" entrytime="00:01:35.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Xenia" lastname="Zolliker" birthdate="2010-10-19" gender="F" nation="SUI" license="7645" swrid="5312756" athleteid="13969">
              <RESULTS>
                <RESULT comment="505 - Wechselbeinschlag während des Schwimmens (Zeit: 8:53)" eventid="1068" status="DSQ" swimtime="00:01:53.43" resultid="13970" heatid="14519" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.51" />
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1078" points="183" swimtime="00:01:36.57" resultid="13971" heatid="14547" lane="2" entrytime="00:01:42.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:36.74" />
                    <SPLIT distance="75" swimtime="00:01:12.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="159" swimtime="00:01:54.97" resultid="13972" heatid="14601" lane="2" entrytime="00:01:59.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:25.17" />
                    <SPLIT distance="50" swimtime="00:00:53.63" />
                    <SPLIT distance="75" swimtime="00:01:25.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="207" swimtime="00:01:24.84" resultid="13973" heatid="14656" lane="1" entrytime="00:01:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.27" />
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="75" swimtime="00:01:03.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="74" swimtime="00:03:14.14" resultid="13974" heatid="14581" lane="2" entrytime="00:02:56.58">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.70" />
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                    <SPLIT distance="75" swimtime="00:01:06.70" />
                    <SPLIT distance="100" swimtime="00:01:30.34" />
                    <SPLIT distance="125" swimtime="00:01:52.10" />
                    <SPLIT distance="150" swimtime="00:02:18.71" />
                    <SPLIT distance="175" swimtime="00:02:44.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13956" number="1" />
                    <RELAYPOSITION athleteid="13952" number="2" />
                    <RELAYPOSITION athleteid="13944" number="3" />
                    <RELAYPOSITION athleteid="13941" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="468" swimtime="00:01:56.44" resultid="13975" heatid="14736" lane="3" entrytime="00:01:58.32">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.34" />
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="75" swimtime="00:00:45.33" />
                    <SPLIT distance="100" swimtime="00:01:02.97" />
                    <SPLIT distance="125" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:31.21" />
                    <SPLIT distance="175" swimtime="00:01:43.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13859" number="1" />
                    <RELAYPOSITION athleteid="13922" number="2" />
                    <RELAYPOSITION athleteid="13931" number="3" />
                    <RELAYPOSITION athleteid="13903" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" points="456" swimtime="00:02:12.96" resultid="13976" heatid="14732" lane="3" entrytime="00:02:15.47">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.43" />
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="75" swimtime="00:00:49.49" />
                    <SPLIT distance="100" swimtime="00:01:09.12" />
                    <SPLIT distance="125" swimtime="00:01:24.88" />
                    <SPLIT distance="150" swimtime="00:01:44.14" />
                    <SPLIT distance="175" swimtime="00:01:57.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13864" number="1" />
                    <RELAYPOSITION athleteid="13936" number="2" />
                    <RELAYPOSITION athleteid="13882" number="3" />
                    <RELAYPOSITION athleteid="13891" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="195" swimtime="00:02:39.28" resultid="13977" heatid="14579" lane="4" entrytime="00:02:43.85">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.19" />
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                    <SPLIT distance="75" swimtime="00:00:56.67" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="125" swimtime="00:01:37.34" />
                    <SPLIT distance="150" swimtime="00:01:59.34" />
                    <SPLIT distance="175" swimtime="00:02:17.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13969" number="1" />
                    <RELAYPOSITION athleteid="13895" number="2" />
                    <RELAYPOSITION athleteid="13914" number="3" />
                    <RELAYPOSITION athleteid="13927" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1084" points="77" swimtime="00:03:36.83" resultid="13978" heatid="14577" lane="2" entrytime="00:02:56.13">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.89" />
                    <SPLIT distance="50" swimtime="00:00:53.57" />
                    <SPLIT distance="75" swimtime="00:01:14.43" />
                    <SPLIT distance="100" swimtime="00:01:43.90" />
                    <SPLIT distance="125" swimtime="00:02:04.15" />
                    <SPLIT distance="150" swimtime="00:02:32.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13869" number="1" />
                    <RELAYPOSITION athleteid="13899" number="2" />
                    <RELAYPOSITION athleteid="13965" number="3" />
                    <RELAYPOSITION athleteid="13851" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Annick" gender="F" lastname="Willemsen" nation="NED" license="7592" />
            <COACH firstname="Agnieszka" gender="F" lastname="Bujoczek" nation="POL" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="STKP" nation="SUI" region="RZW" clubid="13802" swrid="65715" name="Schwimmteam Kaiseraugst-Pratteln" name.en="Stkp" shortname="Stkp">
          <ATHLETES>
            <ATHLETE firstname="Sriraam" lastname="Sivasundaran" birthdate="2007-01-23" gender="M" nation="SUI" swrid="5242675" athleteid="13824">
              <RESULTS>
                <RESULT eventid="1127" points="191" swimtime="00:01:35.95" resultid="13825" heatid="14755" lane="3" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.88" />
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="75" swimtime="00:01:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="208" swimtime="00:01:15.79" resultid="13826" heatid="14785" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.25" />
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="75" swimtime="00:00:55.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Abinaja" lastname="Sivasundaran" birthdate="2008-08-24" gender="F" nation="SUI" swrid="5511492" athleteid="13821">
              <RESULTS>
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="13822" heatid="14706" lane="4" entrytime="00:01:31.00" />
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="13823" heatid="14767" lane="1" entrytime="00:01:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lisa" lastname="Matter" birthdate="2011-01-02" gender="F" nation="SUI" swrid="5085917" athleteid="13807">
              <RESULTS>
                <RESULT eventid="1078" points="167" swimtime="00:01:39.51" resultid="13808" heatid="14548" lane="4" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.93" />
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                    <SPLIT distance="75" swimtime="00:01:14.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="139" swimtime="00:02:00.18" resultid="13809" heatid="14601" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.96" />
                    <SPLIT distance="50" swimtime="00:00:55.52" />
                    <SPLIT distance="75" swimtime="00:01:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="197" swimtime="00:01:26.28" resultid="13810" heatid="14652" lane="4" entrytime="00:01:31.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="75" swimtime="00:01:03.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Weichsel" birthdate="2013-06-06" gender="M" nation="SUI" swrid="5300110" athleteid="13827">
              <RESULTS>
                <RESULT eventid="1100" points="125" swimtime="00:00:40.31" resultid="14510" heatid="14641" lane="3" entrytime="00:00:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="98" swimtime="00:00:48.12" resultid="14511" heatid="14537" lane="3" entrytime="00:00:49.00" />
                <RESULT eventid="1090" points="94" swimtime="00:00:55.34" resultid="14512" heatid="14594" lane="1" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thea" lastname="Richards" birthdate="2010-04-12" gender="F" nation="SUI" swrid="4856317" athleteid="13818">
              <RESULTS>
                <RESULT eventid="1078" points="183" swimtime="00:01:36.55" resultid="13819" heatid="14549" lane="2" entrytime="00:01:36.70">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.90" />
                    <SPLIT distance="50" swimtime="00:00:47.27" />
                    <SPLIT distance="75" swimtime="00:01:12.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="212" swimtime="00:01:24.19" resultid="13820" heatid="14653" lane="2" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.39" />
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                    <SPLIT distance="75" swimtime="00:01:02.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eliza" lastname="Osmani" birthdate="2008-03-05" gender="F" nation="SUI" swrid="5313495" athleteid="13811">
              <RESULTS>
                <RESULT eventid="1114" points="199" swimtime="00:01:33.88" resultid="13812" heatid="14705" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.56" />
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="250" swimtime="00:01:19.73" resultid="13813" heatid="14767" lane="3" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.70" />
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                    <SPLIT distance="75" swimtime="00:00:58.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jasin Tri Thien" lastname="Osmani" birthdate="2010-09-22" gender="M" nation="SUI" swrid="5511488" athleteid="13814">
              <RESULTS>
                <RESULT eventid="1081" points="98" swimtime="00:01:44.52" resultid="13815" heatid="14566" lane="1" entrytime="00:01:49.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                    <SPLIT distance="75" swimtime="00:01:17.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="114" swimtime="00:01:53.87" resultid="13816" heatid="14621" lane="2" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.92" />
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                    <SPLIT distance="75" swimtime="00:01:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="112" swimtime="00:01:33.15" resultid="13817" heatid="14673" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:20.18" />
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                    <SPLIT distance="75" swimtime="00:01:09.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Wüthrich" birthdate="2008-10-22" gender="M" nation="SUI" swrid="5403883" athleteid="13835">
              <RESULTS>
                <RESULT eventid="1111" points="115" swimtime="00:01:37.98" resultid="13836" heatid="14696" lane="1" entrytime="00:01:33.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.10" />
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="75" swimtime="00:01:06.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="230" swimtime="00:01:13.31" resultid="13837" heatid="14787" lane="4" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.52" />
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Weichsel" birthdate="2010-08-31" gender="F" nation="SUI" swrid="4856542" athleteid="13831">
              <RESULTS>
                <RESULT eventid="1078" points="153" swimtime="00:01:42.52" resultid="13832" heatid="14548" lane="1" entrytime="00:01:41.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:23.48" />
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="178" swimtime="00:01:50.81" resultid="13833" heatid="14601" lane="1" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.49" />
                    <SPLIT distance="50" swimtime="00:00:52.49" />
                    <SPLIT distance="75" swimtime="00:01:21.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="197" swimtime="00:01:26.28" resultid="13834" heatid="14653" lane="4" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="75" swimtime="00:01:03.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Demian Alexander" lastname="Dührkop" birthdate="2011-09-24" gender="M" nation="GER" swrid="5223392" athleteid="13803">
              <RESULTS>
                <RESULT eventid="1081" points="117" swimtime="00:01:38.55" resultid="13804" heatid="14565" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.78" />
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                    <SPLIT distance="75" swimtime="00:01:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="78" swimtime="00:02:09.49" resultid="13805" heatid="14619" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.77" />
                    <SPLIT distance="50" swimtime="00:00:56.76" />
                    <SPLIT distance="75" swimtime="00:01:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="105" swimtime="00:01:34.98" resultid="13806" heatid="14676" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.06" />
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="75" swimtime="00:01:08.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Zurflueh" birthdate="2012-10-10" gender="F" nation="SUI" swrid="5403873" athleteid="13838">
              <RESULTS>
                <RESULT eventid="1078" points="170" swimtime="00:01:39.05" resultid="13839" heatid="14549" lane="3" entrytime="00:01:37.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.64" />
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                    <SPLIT distance="75" swimtime="00:01:12.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="157" swimtime="00:01:55.46" resultid="13840" heatid="14602" lane="3" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:24.95" />
                    <SPLIT distance="50" swimtime="00:00:55.89" />
                    <SPLIT distance="75" swimtime="00:01:25.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="193" swimtime="00:01:26.88" resultid="13841" heatid="14652" lane="1" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.53" />
                    <SPLIT distance="50" swimtime="00:00:40.29" />
                    <SPLIT distance="75" swimtime="00:01:03.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="206" swimtime="00:02:36.38" resultid="13842" heatid="14579" lane="2" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.36" />
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                    <SPLIT distance="75" swimtime="00:00:59.08" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="125" swimtime="00:01:37.80" />
                    <SPLIT distance="150" swimtime="00:01:58.54" />
                    <SPLIT distance="175" swimtime="00:02:16.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13838" number="1" />
                    <RELAYPOSITION athleteid="13831" number="2" />
                    <RELAYPOSITION athleteid="13807" number="3" />
                    <RELAYPOSITION athleteid="13818" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4788" nation="GER" region="01" clubid="12852" swrid="67644" name="SSV Grenzach">
          <ATHLETES>
            <ATHLETE firstname="Jan" lastname="Draeger" birthdate="1993-01-01" gender="M" nation="GER" license="135001" swrid="4076925" athleteid="12853">
              <RESULTS>
                <RESULT eventid="1133" points="562" swimtime="00:00:54.45" resultid="12854" heatid="14796" lane="3" entrytime="00:00:54.60">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:11.68" />
                    <SPLIT distance="50" swimtime="00:00:25.19" />
                    <SPLIT distance="75" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="415" swimtime="00:00:29.78" resultid="14856" heatid="14843" lane="1" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Löwe" birthdate="2000-01-01" gender="M" nation="GER" license="322627" swrid="5014453" athleteid="12855">
              <RESULTS>
                <RESULT eventid="1127" points="627" swimtime="00:01:04.63" resultid="12856" heatid="14763" lane="2" entrytime="00:01:03.33">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.59" />
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                    <SPLIT distance="75" swimtime="00:00:46.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="6687" points="343" swimtime="00:00:31.74" resultid="14853" heatid="14802" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="RHYS" nation="SUI" region="ROS" clubid="13176" swrid="65674" name="Rhy Swimming">
          <ATHLETES>
            <ATHLETE firstname="Leonie" lastname="Halter" birthdate="2006-06-07" gender="F" nation="SUI" license="105065" swrid="5073307" athleteid="13186">
              <RESULTS>
                <RESULT eventid="1108" points="318" swimtime="00:01:19.94" resultid="13187" heatid="14687" lane="1" entrytime="00:01:27.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.73" />
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="75" swimtime="00:00:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="410" swimtime="00:01:07.64" resultid="13188" heatid="14775" lane="2" entrytime="00:01:07.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:14.96" />
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="75" swimtime="00:00:50.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andri" lastname="Halter" birthdate="2008-09-19" gender="M" nation="SUI" license="111921" swrid="4821664" athleteid="13183">
              <RESULTS>
                <RESULT eventid="1117" points="338" swimtime="00:01:09.34" resultid="13184" heatid="14726" lane="3" entrytime="00:01:09.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.93" />
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="75" swimtime="00:00:51.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="397" swimtime="00:01:01.10" resultid="13185" heatid="14792" lane="1" entrytime="00:01:01.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.72" />
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                    <SPLIT distance="75" swimtime="00:00:45.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enya" lastname="Buschor" birthdate="2008-10-18" gender="F" nation="SUI" license="112499" swrid="4889092" athleteid="13180">
              <RESULTS>
                <RESULT eventid="1108" status="WDR" swimtime="00:00:00.00" resultid="13181" entrytime="00:01:19.86" entrycourse="SCM" />
                <RESULT eventid="1130" status="WDR" swimtime="00:00:00.00" resultid="13182" entrytime="00:01:09.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Florina" lastname="Wohlgensinger" birthdate="2010-04-09" gender="F" nation="SUI" license="116252" swrid="5261574" athleteid="13195">
              <RESULTS>
                <RESULT eventid="1092" points="380" swimtime="00:01:26.02" resultid="13196" heatid="14610" lane="1" entrytime="00:01:28.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.83" />
                    <SPLIT distance="50" swimtime="00:00:41.17" />
                    <SPLIT distance="75" swimtime="00:01:03.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="307" swimtime="00:01:20.88" resultid="13198" heatid="14522" lane="1" entrytime="00:01:23.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:17.33" />
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="75" swimtime="00:00:59.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="400" swimtime="00:01:08.16" resultid="13199" heatid="14661" lane="1" entrytime="00:01:09.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.66" />
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="75" swimtime="00:00:50.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jasmin" lastname="Weiss" birthdate="2010-08-23" gender="F" nation="GER" license="116248" swrid="5261573" athleteid="13192">
              <RESULTS>
                <RESULT eventid="1092" points="217" swimtime="00:01:43.65" resultid="13193" heatid="14605" lane="4" entrytime="00:01:46.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:21.96" />
                    <SPLIT distance="50" swimtime="00:00:48.17" />
                    <SPLIT distance="75" swimtime="00:01:15.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="247" swimtime="00:01:20.07" resultid="13194" heatid="14658" lane="4" entrytime="00:01:21.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.07" />
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="75" swimtime="00:00:59.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felix" lastname="Weiss" birthdate="2006-07-25" gender="M" nation="SUI" license="101470" swrid="4982697" athleteid="13189">
              <RESULTS>
                <RESULT eventid="1127" points="312" swimtime="00:01:21.55" resultid="13190" heatid="14760" lane="3" entrytime="00:01:21.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.72" />
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                    <SPLIT distance="75" swimtime="00:00:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="393" swimtime="00:01:01.35" resultid="13191" heatid="14792" lane="2" entrytime="00:01:00.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:13.66" />
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="75" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonie" lastname="Billeter" birthdate="2009-11-12" gender="F" nation="SUI" license="111916" swrid="4821662" athleteid="13177">
              <RESULTS>
                <RESULT eventid="1114" points="342" swimtime="00:01:18.43" resultid="13178" heatid="14710" lane="3" entrytime="00:01:20.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:18.52" />
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="75" swimtime="00:00:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="425" swimtime="00:01:06.83" resultid="13179" heatid="14776" lane="2" entrytime="00:01:06.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:15.33" />
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                    <SPLIT distance="75" swimtime="00:00:49.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ladina" lastname="Wohlgensinger" birthdate="2008-02-29" gender="F" nation="SUI" license="111915" swrid="4821671" athleteid="13200">
              <RESULTS>
                <RESULT eventid="1114" points="276" swimtime="00:01:24.27" resultid="13201" heatid="14708" lane="2" entrytime="00:01:23.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:19.27" />
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="75" swimtime="00:01:02.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="262" swimtime="00:01:18.50" resultid="13202" heatid="14769" lane="3" entrytime="00:01:15.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="25" swimtime="00:00:16.52" />
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="75" swimtime="00:00:57.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1120" status="WDR" swimtime="00:00:00.00" resultid="13203" entrytime="00:02:23.68">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13177" number="1" />
                    <RELAYPOSITION athleteid="13186" number="2" />
                    <RELAYPOSITION athleteid="13180" number="3" />
                    <RELAYPOSITION athleteid="13200" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Johanna" gender="F" lastname="Wohlgensinger" type="HEADCOACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="13205" firstname="Billeter" gender="F" lastname="Karin" nation="SUI" />
            <OFFICIAL officialid="13206" firstname="Ladina" gender="F" lastname="Wohlgensinger" nation="SUI" license="111915" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="UNATTACHED">
          <ATHLETES>
            <ATHLETE firstname="Maxime" lastname="Mustermann" birthdate="2007-01-01" gender="F" athleteid="14490">
              <RESULTS>
                <RESULT eventid="6681" swimtime="00:00:00.00" resultid="14492" entrytime="00:02:30.00" />
                <RESULT eventid="6635" swimtime="00:00:00.00" resultid="14493" entrytime="00:02:30.00" />
                <RESULT eventid="6637" swimtime="00:00:00.00" resultid="14494" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Max" lastname="Mustermann" birthdate="2007-01-01" gender="M" athleteid="14489">
              <RESULTS>
                <RESULT eventid="6687" status="DNS" swimtime="00:00:00.00" resultid="14495" entrytime="00:02:30.00" />
                <RESULT eventid="6683" swimtime="00:00:00.00" resultid="14496" entrytime="00:02:30.00" />
                <RESULT eventid="6639" swimtime="00:00:00.00" resultid="14497" entrytime="00:02:30.00" />
                <RESULT eventid="6679" swimtime="00:00:00.00" resultid="14498" entrytime="00:02:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maxime" lastname="Mustermann" birthdate="2010-01-01" gender="F" athleteid="14500" />
            <ATHLETE firstname="Max" lastname="Mustermann" birthdate="2010-01-01" gender="M" athleteid="14499" />
          </ATHLETES>
          <OFFICIALS>
            <OFFICIAL officialid="14834" firstname="Francesca" gender="F" lastname="Garotta" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
